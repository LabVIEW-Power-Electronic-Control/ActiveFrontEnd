-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��b�d�l��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e��!�:�$�8�G��6����g"��x)��*�����}�d�3�*����P���F��1�����&�0�e�4��1�W���,�Ɵ�w9��p'�����u�
�
�6�>�3�(���Y�ƃ�gF��s1��2������u�d�}�������9F���*���<�;�
�
��-����Cө��5��h"��<��u�u�%�e��)�������)��=��*����
����u�FϺ�����O��N������!�:�&�2�o��������|3��d:��9����_�u�u���������� F��x;��&���������W��Y����G	�UךU���
�
�6�<�9��(܁�	����\��b:��!�����n�u�w�-�G�������l��T�� ����
�����#���Q����\��XN�N���u�%�e��#�2����M����E
��N��!ʆ�����]�}�W���&����\��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
��>����&����R��[
��U���u��
���f�W���	�֓�P��Y��*���u� �u����>���<����N��
�����e�n�u�u�'�m�6�������lP��G1����������4�ԜY�Ƽ�9��C�����b�o�����;���:����g)��]����!�u�|�_�w�}�(߁�����@9�� 1��*���u�u� �u���8���B�����h/�����
�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�I����Z	��h��*���#�1�o����3���>����F�G1��4���:�&�0�l�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����r��X �����4�
�9�u�w��W���&����p]ǻN��*ي� �%�!�
��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lU��B�����
�
�%�#�3�g�8���*����|!��d��Uʥ�f��!� �$�8�F��6����g"��x)��*�����}�d�3�*����P���F��1�����&�0�d�4��1�W���,�Ɵ�w9��p'�����u�
�
� �'�)�(���Y�ƃ�gF��s1��2������u�d�}�������9F���*���%�!�
�
��-����Cө��5��h"��<��u�u�%�f��)�������)��=��*����
����u�FϺ�����O��N������!� �&�2�n��������|3��d:��9����_�u�u����������F��x;��&���������W��Y����G	�UךU���
�
� �%�#��(ہ�	����\��b:��!�����n�u�w�-�D�������l��T�� ����
�����#���Q����\��XN�N���u�%�f��#�(����L����E
��N��!ʆ�����]�}�W���&����F��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
��(����&����R��[
��U���u��
���f�W���	�Փ�F��C��*���u� �u����>���<����N��
�����e�n�u�u�'�n�8�������lQ��G1����������4�ԜY�Ƽ� 9��C�����m�o�����;���:����g)��]����!�u�|�_�w�}�(܁�����@9��1��*���u�u� �u���8���B�����h!�����
�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�J����C��h��*���#�1�o����3���>����F�G1��:��� �&�0�d�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l)��G��*���e�4�
�9�w�}�"���-����t/��=N��U���
�4� �9�8�)����&����z(��c*��:���n�u�u�4��8�Mϗ�Y����)��tUךU���
�
�4� �;�2����&����R��[
��U��������W�W���&ǹ��]��t�����0�d�o��w�	�(���0����p2��F�U���;�:�e�n�w�}����4����_%��C��*���
�%�#�1�m��W���&����p]ǻN��*ފ�4� �9�:�#�2�(���Y�ƅ�5��h"��<��u�u�%�a��3��������l��h�����o��u����>��Y����lR��V �����!�:�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����~��V�����9�0�f�4��1�W���7ӵ��l*��~-�U���%�a��;�6���������\��yN��1�����_�u�w��(�������]��[1��A���
�9�u�u���3���>����F�G1��8���4��;�'�;�8�B��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����h#�� ���:�!�:�
����������}F��s1��2���_�u�u�
��<��������_9��N�<����
���l�}�WϮ�M����F��X �����
�
�%�#�3�g�>���-����t/��=N��U���
�4� �9�8�)����&����z(��c*��:���
�����l��������l�N��A���;�4��;�%�1��������WF��~ ��!�����n�u�w�-�B�������lV�'��&���������W��Y����G	�UךU���
�
�4�2���(������/��d:��9����_�u�u������&����	F��=��*����
����u�FϺ�����O��N������;�0�0�f�<�(���Y�ƅ�5��h"��<��u�u�%�`��3����K����}F��s1��2������u�d�}�������9F���*���2�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�4�0��(���Y����g"��x)��*�����}�d�3�*����P���F��1�����0�f�4�
�;�}�W���*����|!��d��Uʥ�`��;�0�2�i�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����lS��V ��*���
�%�#�1�m��W���&����p]ǻN��*ߊ�4�2�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����a��R1��@���
�9�u�u���3���>����F�G1��'���0�0�c�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�L����T��hX�����1�o��u���8���B�����h<�����
�u�u����;���:����g)��]����!�u�|�_�w�}�(ځ�����V9��V�����u������4�ԜY�Ƽ�9��Y	����o��u����>���<����N��
�����e�n�u�u�'�h�%�������l��A��Oʜ�u��
���f�W���	�ӓ�R��h��U���������!���6���F��@ ��U���_�u�u�
��<����&ʹ��l��T��;ʆ�����]�}�W���&����^��E��*���u������4���:����U��S�����|�_�u�u����������l��h�����o��u����>��Y����lP��V�����&�0�d�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�O����R��R�����4�
�9�u�w��$���5����l�N��C���'�8�!�'���W���7ӵ��l*��~-��0����}�u�:�9�2�G��Y����lP��V�����&�0�g�4��1�W���7ӵ��l*��~-�U���%�c��'�:�)����&����z(��c*��:���
�����}�������9F���*���4�0�0�&�2�n��������z(��c*��:���n�u�u�%�`��������/��d:��9�������w�n�W������]ǻN��*݊�4�;�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�
�6�3�(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�G1��2���&�0�d�4��1�W���7ӵ��l*��~-�U���%�b��<�$�8�E��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����h)�����
�
�%�#�3�g�>���-����t/��=N��U���
�4�;�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�Ƽ�9��^ �����4�
�9�u�w��$���5����l�N��B���<�&�0�a�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ѓ�R��h��*���#�1�o��w�	�(���0��ƹF��hY�����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����@9��1��*���u�u�����0���s���C9��p�����c�o��u���8���&����|4�_�����:�e�n�u�w�-�@�������lP��G1�����u��
���L���YӖ��l!��Y��*���u������4���:����U��S�����|�_�u�u������&����R��[
��U��������W�W���&Ĺ��Z��R1�Oʜ�u��
����2���+������Y��E��u�u�%�b��4����A����E
��N��U���
���n�w�}����>����l��T��;ʆ�������8���J�ƨ�D��^����u�
�
�4�9��(ց�	����\��yN��1�����_�u�w��(�������V9��N��U���
���n�w�}����*����_��h^�����1�o��u���8���B�����h=�����
�
�u�u���3���>����F�G1��&���4�&�0�d�6�����Y����g"��x)��N���u�%�d�
�2�-����&����	F��=��*����
����u�FϺ�����O��N����
�0�%�<�#��(߁�	����\��yN��1�����_�u�w��G�������G��h_��U���������4���Y����W	��C��\�ߊu�u�
�e��)����
����l��A��Oʜ�u��
���f�W���	����z��C��*���u������4���:����U��S�����|�_�u�u��l�>�������9��h��U���������}���Y����l/��B����o��u����>���<����N��
�����e�n�u�u�'�l�(�������lW��G1�����u��
���L���YӖ��9��G��*���u�u�����0���/����aF�N�����u�|�_�u�w��F���	����V9��V�����u������4�ԜY�Ƽ�W��Y�����f�o��u���8���&����|4�_�����:�e�n�u�w�-�Fށ�����l��h�����o��u����>��Y����lW��~ �����
�u�u����;���:����g)��]����!�u�|�_�w�}�(���0����@9��1��*���u�u�����0���s���C9��h'�� ���0�`�o��w�	�(���0����p2��F�U���;�:�e�n�w�}���&����G��h[�����1�o��u���8���B�����1�����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���H����F��R1�����9�u�u����;���:����V��=d�����!�6� �0�5�5�ϱ�Y�֍�S����U���_�u�u�!�%�?����6����v(��v:��;����u�u����}���Y����Z��RN��'���������1���ӄ��R������6� �0�<�]�}�Wͳ�8����_��B�����
�e�a�a�,��(���,����c#��O��9���� �
���`�[���&����g9��o+��EƝ�������J�������_��C�=���������E���I����.��h'�� �����:�=�%�q�;��� ����|%��_�E��e������#��J߮��l5��h:��H���0������:��U����`?��s=��F����
��
��k�N���5����}9��cS�B���w�_�u�u�8�.��������]��[����o������M���H��ƹF��X �����4�
�:�&��2����Y�Ɵ�w9��p'��O���e�n�u�u�4�3����Y����g9��1����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-�$�������^9��N��1��������}�E�������V�S��E��e�e�e�e�g�m�G��H����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�g�u�8�3���Y���V��^�E��e�e�e�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�w�_�u�w�2����Ӈ��`2��C[�����u�u��
���(���-���W��X����u�h�w�e�g�m�G��I����W��^�����u�:�&�4�#�<�(���
�Г�@��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I���9F������!�4�
��$�j����O����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�d�e�g�m�L���YӅ��@��CN��*���&�m�3�8�`�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�����m�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�N���u�6�;�!�9�}����&����l ��hW��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
��.�Fށ�
����\��c*��:���
�����l��������\�^�E��e�e�d�e�g�m�G��B�����D��ʴ�
��&�d��.�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�f�W�������R��V��!���d�
�&�
�e�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�*���
�f�o����0���/����aF�N�����u�|�o�u�g�m�G��H����V��^�E��u�u�6�;�#�3�W���*����S��D��A��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'��(���O����lW��N��1��������}�E�������V�S��E��e�d�e�e�g�m�G��I����F�T�����u�%��
�#�j����H����`2��{!��6�����u�g�w�2����I����D��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�m�3�:�l�W���-����t/��a+��:���g�u�:�;�8�m�W��[����V��^�E��e�e�e�w�]�}�W���
������d:�����3�8�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��w�_�u�u�8�.��������l��1����u�u��
���(���-���W��X����u�h�w�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����U��^��U���
���
��	�%���Hӂ��]��G��H���d�e�e�e�g�m�G��I����]ǻN�����4�!�4�
��.�E݁�
����\��c*��:���
�����l��������\�_�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�G��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�e�1�"�#�}�^��Y���9F������!�4�
�:�$�����J����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lQ�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��_�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h+��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��\��G��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��e�n�u�u�4�3����Y����\��h��G��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�d�n�u�w�>�����ƭ�l��D������o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��X ��*���g��o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�d�d�l�}�WϽ�����GF��h�����#�g�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�f�
�d�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�m�F��Y����\��V �����:�&�
�#�e��Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�F��B�����D��ʴ�
�:�&�
�!�o�F���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>��������  ��t*�U����
�����#���Q����\��XN�U��w�e�d�d�f�m�F��H����W��^�E��w�_�u�u�8�.��������]��[�*ٓ��a�e�o���;���:����g)��]����!�u�|�o�w�m�F��H����W��_�D��e�e�e�e�g�f�W�������R��V�����
�#�g�f���6���Y����)��t1��6���u�f�u�:�9�2�G���D����W��^�D��d�d�d�d�f�l�F��H����F�T�����u�%�6�;�#�1�D݁�N����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��H����]ǻN�����4�!�4�
�8�.�(���K�׉�	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>�����ޓ�\��c*��:���
�����}�������	[�^�E��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��^��U���
���
��	�%���Mӂ��]��G��H���e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�f��C��Cӵ��l*��~-��0����}�a�1� �)�W���C���V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��M���u�u��
���(���-���F��@ ��U���o�u�d�d�f�l�U�ԜY�Ư�]��Y�����;�!�9�d��m�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��n�u�u�6�9�)����	����@��A_��D��o������!���6���F��@ ��U���o�u�e�e�g�l�G��I���9F������!�4�
�:�$�����M���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����d�
�u�u���8���&����|4�N�����u�|�o�u�g�m�G��I����F�T�����u�%�6�;�#�1�Fׁ�Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�e�w�]�}�W���
������T�����d�
��o���;���:����g)��_����!�u�|�o�w�m�G��I����W��_�N���u�6�;�!�9�}��������EW��(��3��������4���Y����W	��C��\��u�d�d�d�f�l�F��H����l�N�����;�u�%�6�9�)���&����V��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W��n�u�u�6�9�)����	����@��A\��U����
�����#���Q�ƨ�D��^��O���e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}�����ƭ�l%��Q��Oʆ�������8���K�ƨ�D��^��O���e�e�e�e�g�m�G��I����D��N�����<� �0�3�:�8��������@��Y	�U���4�!�<� �2�;��������TF����6���&�u�u�<�9�1��������l�N�����u�%�&�2�4�8�(���
�ד�@��T��!�����n�u�w�.����Y����Z��S
��M������]�}�W�������lR��V �����!�:�
�
��3����Cӵ��l*��~-�U���&�2�4�u����������A	��R1�����u�u��
���W��^����F�D�����
�
�4� �;�2����&����R��[
�����2�o�����4�ԜY�ƿ�T����*��� �9�:�!�8��(߁�	����l��PN�&������o�w�m�L���Yӕ��]��G1��8���4��;�'�;�8�F���&����	F��s1��2������u�d�}�������9F������%�a��;�6���������l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�&�2�6�}�(ہ�����p	��E�����4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
��<��������_9��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�a��3��������l��h�����o������}���Y����R
��hZ�����9�:�!�:���(�������g"��x)��U��r�r�_�u�w�4����	�ғ�R��[-�����
�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�C�������\��X��*؊�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��(�������]��[1��F���
�<�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����~��V�����9�0�f�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*ފ�4� �9�:�#�2�(���&����_��Y1���������W�W���������h#�� ���:�!�:�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��z�����;�'�9�0�c�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�i�:�������G��h��*���2�o�����4��Y���9F������%�a��;�6���������l��A�����<�u�u����>��Y����Z��[N��A���;�4��;�%�1��������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*��� �9�:�!�8��(ځ�����\��c*��:���
�����l��������l�N�����u�
�
�4�"�1��������9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1����4����_%��C��*���
�%�#�1�>�����Y����)��tUךU���<�;�9�%�c�����:����\
��h[�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��<��������_9��1��*���u�u��
���L���Yӕ��]��G1��8���4��;�'�;�8�A�������`2��{!��6��u�e�n�u�w�.����Y����~��V�����9�0�c�4��1�(���
���5��h"��<��u�u�&�2�6�}�(ہ�����p	��E�����4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�C�������\��X��*݊�;�&�2�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l+��B�����:�
�
�
�%�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����Y������;�4��9�/����N����E
��^ �����u��
���f�W���
����_F��1������;�'�9�2�j��������V�=��*����u�h�r�p�W�W���������h<�����
�
�;�&�0�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h<�����
�
�'�2�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�L���Yӕ��]��G1��'���0�0�e�4��1�(���
���5��h"��<��u�u�&�2�6�}�(ځ�����V9��V�����'�2�o����0���C���]ǻN�����9�%�`��9�8��������TF��d:��9�������w�n�W������]ǻN�����9�%�`��9�8����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
��<����&¹��l��h�����o������}���Y����R
��h[�����
�
�
�%�!�9����Y�Ɵ�w9��p'��O���e�n�u�u�$�:����&ƹ��]��R1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ƹ��]��R1�����u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}����Ӗ��l4��P��*؊�%�#�1�<��4�W���-����t/��=N��U���;�9�%�`��3����K����E
��G��U����
���w�`�P���s���@��V��*ߊ�4�2�
�
��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ߊ�4�2�
�
��/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʥ�`��;�0�2�n��������l��T��!�����n�u�w�.����Y����a��R1��F���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�h�%�������l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�h�%�������l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�&�2�6�}�(ځ�����V9��V�����;�&�2�o���;���:���F��P ��U���
�4�2�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��e�����`�<�
�<�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��e�����`�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����R
��h[�����
�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�B�������lS��G1�����0�u�u����>���D����l�N�����u�
�
�4�0��(ف�����\��c*��:���
�����l��������l�N�����u�
�
�4�0��(ف����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�`��3����O����E
��^ �����u��
���f�W���
����_F��1�����0�c�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�L����T��hY�����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�L����T��hY�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����a��R1��B���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�6�:�(���&����_��E��Oʆ�����m�}�G��Y����Z��[N��@���;�0�0�m�>�����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��@���;�0�0�m�'�8�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��P ��U���
�4�2�
����������@��N��1�����_�u�w�4����	�ӓ�R��h��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u������&����Z��^	��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u������&����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�<�;�;�-�B�������l_��G1�����
�<�u�u���8���B�����Y������;�0�0�n�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lP��V�����&�0�e�<��4�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��%���8�!�'�
������Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������%�c��'�:�)����&ù��l��h�����o������}���Y����R
��hX�����0�0�&�0�g�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lP��V�����&�0�d�<��4�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��%���8�!�'�
������Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������%�c��'�:�)����&¹��l��h�����o������}���Y����R
��hX�����0�0�&�0�f�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lQ��V��*���
�;�&�2�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������lQ��V��*���
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F�� 1�����0�e�4�
�;���������g"��x)��N���u�&�2�4�w��(�������9��h��*���2�o�����4��Y���9F������%�b��<�$�8�F���&����	F��s1��2������u�d�}�������9F������%�b��<�$�8�F�������`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����4�u�
�
�6�3�(���&����_��Y1���������W�W���������h)�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����@9��1��*���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����@9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ѓ�R��h��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�b��>�.��������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*���;�
�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���;�
�
�
�%�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����Y������<�&�0�d�<�(���&����Z�=��*����n�u�u�$�:����&Ĺ��Z��R1�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�`������ғ�]9��PN�&���������W��Y����G	�UךU���<�;�9�%�`������ғ�A��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�&�2�4�w��(�������9��h��*���&�2�o����0���s���@��V��*݊�4�;�
�
��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��^ �����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��^ �����%�0�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W���������h)�����
�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�j�0���
����l��A�����u�u��
���W��^����F�D�����
�
�4�;���(���
���5��h"��<������}�f�9� ���Y����F�D�����
�
�4�;���(�������g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����9�%�b��>�.��������W9��h��U����
���l�}�Wϭ�����C9��p�����c�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����>����l��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����>����l��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:����&Ĺ��Z��R1�����9�
�;�&�0�g�$���5����l�N�����u�
�
�4�9��(؁�	����l��PN�&������o�w�m�L���Yӕ��]��G1��2���&�0�m�<��4�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��2���&�0�m�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*݊�4�;�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�N����]��hV�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��<����&ʹ��l��T��!�����
����_������\F��d��Uʦ�2�4�u�
��<����&ʹ��V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�<�;�9�'�j�0���
����l��A�����<�u�u����>��Y����Z��[N��B���<�&�0�l�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l5��Y��*���
�;�&�2�m��3���>����F�D�����
�
�<�;�;��(߁����5��h"��<���h�r�r�_�w�}����Ӗ��l5��Y��*���
�%�#�1�>�����Y����)��tUךU���<�;�9�%�n�����
����l��A�����u�u��
���W��^����F�D�����
�
�<�;�;��(ށ�����\��c*��:���n�u�u�&�0�<�W���&����R
��R1�����u�u��
���W��^����F�D�����
�
�<�;�;��(ށ�	����l��D��Oʆ�����]�}�W�������l_��^	�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���I����C	��C��*ڊ�;�&�2�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��9��C�����0�e�%�0�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�ƿ�T����E���!�:�;�&�2�m��������l��T��!�����n�u�w�.����Y����l5��G�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���H����F��R1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&�ד�]��D1��E���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W�������lW��~ �����
�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�l�(�������lV��G1�����0�u�u����>���D����l�N�����u�
�d��'�)�(���&����Z�=��*����
����u�FϺ�����O��N�����4�u�
�d��-����&¹��V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�<�;�9�'�l�(�������lW��G1�����
�<�u�u���8���B�����Y����
�;� �&�2�l��������V�=��*����u�h�r�p�W�W���������1�����
�
�
�;�$�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h_��<���!�
�
�
�%�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����Y����
�;� �&�2�o��������l��T��!�����n�u�w�.����Y����l/��B�����4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�Fށ�����l��h�����o������!���6���F��@ ��U���_�u�u�<�9�1���&����G��h]�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����l/��B�����4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
�f�����&����R��[
�����o������M���I��ƹF��^	��ʥ�d�
�;� �$�8�C���&����	F��s1��2������u�d�}�������9F������%�d�
�;�"�.����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
�f�����&����R��[
�����2�o�����4�ԜY�ƿ�T����D���%�!�
�
��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�W��Y�����`�<�
�<�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��h'�� ���0�`�%�0�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�ƿ�T����D���%�!�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�H¹��C��h��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u��l�>�������9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��F���	����V9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�>�3�Ϯ�H¹��C��h��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�d�
�9�(����O����E
��G��U����
���w�`�P���s���@��V��������:�#�(�(���I����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���<�;�9�2�'�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����0�
�g�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�l��h�����
�!�
�&��}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(�������@��Q��C�������W�W���������D�����a�b�o����9�ԜY�ƿ�T�������6�0�
��$�l�(���&���5��h"��<��u�u�&�2�6�}��������lS��T��:����n�u�u�$�:��������lP��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�%�:�@��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V����� �b�b�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����A�� Z�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�����
����g9��1����o������}���Y����R
��G1�����1�`�l�o���2���s���@��V�����
�
�
�e�1��@ׁ�	����VF��d:��9����_�u�u�>�3�Ͽ�&����P��h=�����3�8�m�o���;���:���F��P ��U���&�2�7�1�b�l�MϜ�6����l�N�����u�%�&�2�4�8�(���
����U��Z��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��G1��E���f�3�
�d��-����Y�Ɵ�w9��p'�����u�<�;�9�6�����
����g9��W�����m�o�����4�ԜY�ƿ�T�������7�1�`�f�m��8���7���F��P ��U���
� �b�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��P1�E��������4���Y����W	��C��\�ߊu�u�<�;�;�:����&����CT�=��*����
����u�FϺ�����O��N�����4�u�0�
�b�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������T�=��*����
����u�FϺ�����O��N�����4�u�0�
�a�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��*���$��
�!�g�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������B9��h��D���8�d�u�u���8���B�����Y�����<�
�1�
�`�}�W���5����9F������'�2�b�a�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1����c�o�����}���Y����R
��d1�� ���;� �
�e�f�;�(��&���5��h"��<������}�f�9� ���Y����F�D������-� ��9�(�(���H����lW��N�&���������W��Y����G	�UךU���<�;�9�3���;���6����9��Q��D���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����2��x��Gڊ�
�0�
�c�c�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������q+��7���:�!� �
�`�8�G�������
F��d:��9�������w�n�W������]ǻN�����9�2�%�3��d�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&��� �,� �
�f�l����H����	F��s1��2������u�d�}�������9F������2�%�3�
�n��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������,� �
�f�f�/���O����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
�:�0�!�%�����
����Z9��h��*��c�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����l��Z1�������<�d��8�(��K����g"��x)��*�����}�d�3�*����P���F��P ��U���-� ���#���������9��P1�B���u��
����2���+������Y��E��u�u�&�2�6�}�$���,����F��B�����d�
�
�0��k�D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������,� �
�d�f�/���A����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���M����lW��N��1�����_�u�w�4��������T9��S1�C������]�}�W�������A��h^��*���3�
�c�
�'�9����Y����)��tUךU���<�;�9�3���5�������G��C1�*ۊ�0�
�c�a�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������_9��S������'�0�=�$��;����ד�V�� ^�Oʆ�������8���J�ƨ�D��^����u�<�;�9�4���������g��R>������&�6�g�%�:�F��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����:�0�!�'��5��������9��T1����d�u�u����>���<����N��
�����e�n�u�u�$�:��������V9��E�����1�1�:�!�8��(���&����\��c*��:���
�����l��������l�N�����u�9�;�1��8����
����W%��C��*���
�0�
�b�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������Y��*���8��&�4�2���������l��h_�C��������4���Y����W	��C��\�ߊu�u�<�;�;�>�(�������^9��D�����;�'�9�&�d�/���J����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʶ�
�:�0�!�%���������]��[1��A���2�d�f�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ư�l��R1�����4�6�1�1�8�)����&ƹ��T9��_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�;�3��������R��S�����:�
�
�
�2��@��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����1�
�0�8��.����:����\
��hY�����b�d�o����0���/����aF�N�����u�|�_�u�w�4��������f$��B��*���
�b�c�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�d�
�&��j�Mύ�=����z%��N�����4�u�%�&�0�?���K����|)��v �U���&�2�4�u��%�3�������A��Y�U����
�����#���Q����\��XN�N���u�&�2�4�w�����-����G9��1��*��g�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����~3�� �����d�'�2�d�`�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h �����
�e�3�
�c�d����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�G�������	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������lV��h]�� ��m�4�
�!�%�}�W���&����p]ǻN�����9�2�%�3�g�;�D���&����R��S��Oʆ�����]�}�W�������A��h^��*ي� �c�m�4��8����Y����)��tUךU���<�;�9�2�'�;�G���J����W��^ �����
�
�
�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��1��F���
�d�
�;��3�������5��h"��<������}�f�9� ���Y����F�D�����'�
�
�
�����A����a��R1����o������!���6���F��@ ��U���_�u�u�<�9�1�����֓�lU��B1�M���
�4�2�
���W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�f�3�
�f���������l��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���&����^��Y1�����b�0�`�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��h��*���c�m�<�
�6�:�(؁�&����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�e�3�d�;�(��&����R��hY��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù�� 9��hX�*����;�4��9�/���&����	F��s1��2���_�u�u�<�9�1�����֓�lU��B1�M���
�4� �9�8�)����K����\��c*��:���
�����l��������l�N�����u�'�
�
���(���O�ޓ�]9��Y��6���'�9�d�
��}�W���&����p]ǻN�����9�2�%�3�g�;�D���&����Z��V �����!�:�
�g�2�n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �c�o�4�(�������]��[1�*���u�u��
���L���Yӕ��]��P�����3�f�3�
�f���������\��X��G���`�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����l ��h��C���<�
�4� �;�2����&�ԓ�lP�=��*����n�u�u�$�:��������9��1��*��
�;��;�6���������V9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������9��h)�����
�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����d�
�;��>�.�C���H����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�A�������Z��1��G��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����l ��_�����4�;�
�
��}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���f�3�
�d��3�0���
�ғ�lR�=��*����
����u�FϺ�����O��N�����4�u�'�
���(܁�����l��p�����0�`�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h]�� ��m�<�
�4�9��(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�e�3�f�1��Fׁ�����]��h��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����U��V�����&�!�e�o���;���:���F��P ��U���
�
�
�
��(�A�������lT��h^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��(߁�&����lP��h��%���
�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����d�
�;����(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�f�3��l�(���)����V9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������9��h=��D���e�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����l ��h��C���<�
��d�2�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �c�o�<�(�������\��c*��:���
�����l��������l�N�����u�'�
�
���(���O�ޓ�C9��C��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù�� 9��hX�*���'�!�'�
�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q1�����3�
�d�
�'�/����&����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�e�3�d�;�(��&����V��Y1�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-�����Փ�F9��1��*��� �;�`�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��h��*���c�m�4�
�2�(���Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
�
�
�"�k�O���&����A��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���&����^��G1�����
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�%�'�!�%��W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�f�3�
�f�����Y�Ɵ�w9��p'�����u�<�;�9�0�-��������U��_�����4�!�o����0���s���@��V�����
�
�
�d�1��Aށ�	����VF��d:��9����_�u�u�>�3�Ϲ�	����l ��1��*��
�%�'�4�.�g�$���5����l�N�����u�'�
�
���F���&����Z��{"�����l�0�e�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��h��D���
�c�
�;������&ʹ��F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�Fށ�����l��E����o������}���Y����R
��E��*ڊ�
�d�3�
�a�����5����@9��R1�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-��������U��_������4�;�
���W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�d�
� �a�l��������]9��R1�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-��������U��_�����<��%�6�2�����L����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
�f�;�(��&����g9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m���&����W��Y1��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù��W��B1�D���
�0� �;�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���d�3�
�c��-��������	F��s1��2������u�d�}�������9F������2�%�3�e�1�l�(���O�ד�C9��C��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù��W��B1�D���
�0� �;�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���d�3�
�c��-����Y����)��tUךU���<�;�9�4��4�(�������@��h��*��o������}���Y����R
��G1�����1�m�d�o���2���s���@��V�����
�
�
�e�1��@ׁ�	����A�=��*����n�u�u�$�:��������9��^�� ��m�4�
�1�2�g�$���5����l�N�����u�'�
�
���G���&����R��R��U����
���l�}�Wϭ�����T��Q1����
� �c�m�>��(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�d�
�"�k�O���&����A��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���I����Q��V�����;�d�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h_�����b�
�%�6�w�}�#���6����9F������2�%�3�e�1�n����H˹��l��E�����4�!�'�2�m��3���>���F�UךU���<�;�9�2�'�;�G���H¹��lP��h�����!�4�
�!�%�����Y����)��tN�U��n�u�u�&�0�<�W���&����U9��h��C���4�
�!�'��-��������\��c*��:���u�h�r�r�]�}�W�������C9��P1������&�g�
�$��F��*����|!��d��Uʦ�2�4�u�%�$�:����H����	F��x"��;�ߊu�u�<�;�;�:����&����CV�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�k�@���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����<�
�&�$���݁�
����	F��s1��2���_�u�u�<�9�1��������W9��Y��U�����n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��G��CӤ��#��d��Uʦ�2�4�u�%�$�:����&����GW��Q��D���u��
���f�W���
����_F��h��*���
�e�d�o���2���s���@��V����� �c�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q��Lۊ�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����_��G^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%����L����	F��s1��2������u�d�}�������9F������2�%�3�
�n��G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���c�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��hY�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��(�@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�
�d��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�� ��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U��Y��D��������4���Y����W	��C��\�ߊu�u�<�;�;�:����&����CV�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�j�F���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�
� �`�l����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����3�
�m�
�c�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����_	��a1�*���b�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��^1��Fӊ� �m�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��h��*���b�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӕ��l��h�� ��d�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����U��^1�����
�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G_��*���m�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1�����a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����9��^1�����
�4�!�3��o�(��Cӵ��l*��~-��0����}�a�1� �)�W���s���@��V�����8�
�
� �o�n����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��'���9�
�b�3��k�(��Cӵ��l*��~-��0����}�b�1� �)�W���s���@��V��&��� ��;� ��m��������9��hV�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�l�G�������9��T��!�����
����_�������V�=N��U���;�9�!�%�1��O؁�K����g"��x)��*�����}�u�8�3���B�����Y�����c�
� �l�f�-�W���-����t/��a+��:���b�1�"�!�w�t�}���Y����R
��Z��E؊� �l�l�%�w�}�#���6����e#��x<��Bʱ�"�!�u�|�]�}�W�������^��1��*��
�f�o����0���/����aF�
�����e�n�u�u�$�:����&����lW��h��M���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l��B1�D���u�u��
���(���-��� V��X����n�u�u�&�0�<�W�������l^��Q��Gӊ�`�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����gT��B��E���
�%�,�0�1��B܁�J����g"��x)��*�����}�a�3�*����P���F��P ��U���
�8�c�<�1��Cځ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�
�"�d�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�m�<�3��h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*����g��!�e����H����	F��s1��2������u�d�}�������9F������%��9�
�n�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����:�
�
�e�1��@ځ�M����g"��x)��*�����}�u�8�3���B�����Y������g�
� �n�h����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����<�<�
� �n�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���
�`�3�
�o��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��E�����<�
� �d�g��D��*����|!��h8��!���}�a�1�"�#�}�^�ԜY�ƿ�T����*��
�
�
�m�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�d�<��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�
�c�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����0�
�
�
��d����&����l ��^�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������9��h_�F���u�u��
���(���-���R��X����n�u�u�&�0�<�W�������l^��Q��E���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����2��x��Gڊ�;�0�%��d�;�(��@����	F��s1��2������u�f�}�������9F������!�%�<�
�"�l�Aځ�K����g"��x)��*�����}�u�8�3���B�����Y�����d�e�<�
�"�l�@ށ�K����g"��x)��*�����}�u�8�3���B�����Y�����m�
� �d�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Cފ� �d�l�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��^�����e�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��l^��Q��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�I����9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	����F
��^�� ��d�
�`�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��K+��c\�� ���e�<�
�%�.�8�F���&����l��N��1��������}�F�������V�=N��U���;�9�&�9�#�-�(������� S��N�&���������W������\F��d��Uʦ�2�4�u�0��0�@���&����R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)�ׁ�H����W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��%�"�������V��h��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4����	����9��h��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������lT��Q��G���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϲ����� 9��h_�A���u�u��
���(���-���T��X����n�u�u�&�0�<�W���&����ZW��1��*��a�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l��1��*��m�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l��1��*��e�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����U��^1��ۊ� �d�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���3�
�f�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��G���
� �d�e��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��C1�����<�d�6�&��<����&����l��N��1��������}�F�������V�=N��U���;�9�&�9�#�-�ځ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�2�(��������V��N�&���������W��Y����G	�UךU���<�;�9�3���;���6����l��R��#���3�
�f�m�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��*���d�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1�����f�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��l^��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���O����U��h�Oʆ�������8���Nӂ��]��G�U���&�2�4�u�:��B���&����l��N��1��������}�@Ϻ�����O��N�����4�u�
�g�g�l�݁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��j����&����l��N��1��������}�D�������V�=N��U���;�9�%��$�1�(�������^��N�&���������W��Y����G	�UךU���<�;�9�3���;���6����l��Q����� �d�d�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��C���
� �d�e��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1��݊�g�3�
�a�g�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����<�
� �d�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Q=��8���g��!�b�1��C���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
��-� ��m��������U��\�����u��
����2���+������Y��E��u�u�&�2�6�}�$���>����lW��Y�����
�a�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q��M݊�%�:�0�o���;���:����g)��_�����:�e�n�u�w�.����Y����U��Y���������W�W���������D�����
��&�c�1�0�B��*����|!��d��Uʦ�2�4�u�%�$�:����H����	F��x"��;�ߊu�u�<�;�;�:����&����\��S��U���
���
��	�%���Y����G	�UךU���<�;�9�2�'�;�(��&���5��h"��<��u�u�&�2�6�}��������l��N��1�����_�u�w�4��������F9��1��U����
���l�}�Wϭ�����R��d1����������4���Y����W	��C��\�ߊu�u�<�;�;�<�(���&����V��N��:����_�u�u�>�3�Ͽ�&����Q��\�Oʗ����_�w�}����Ӈ��@��U
��A��o�����W�W���������D�����a�d�o����9�ԜY�ƿ�T�������7�1�a�e�m��8���7���F��P ��U���&�2�7�1�c�d�MϜ�6����l�N�����u�%�&�2�5�9�C��CӤ��#��d��Uʦ�2�4�u�%�$�:����M���$��{+��N���u�&�2�4�w�-��������F��u!��0���_�u�u�<�9�1��������W9�� N�7�����_�u�w�4��������T9��S1�C������]�}�W�������C9��P1����`�o�����}���Y����R
��G1�����1�d�a�o���2���s���@��V�����2�7�1�d�d�g�5���<����F�D�����%�&�2�7�3�l�E��;����r(��N�����4�u�%�&�0�?���H����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:����	����l��h_�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�e�u�u���6��Y����Z��[N��*���
�1�
�d�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����S��N��:����_�u�u�>�3�Ͽ�&����Q��X�Oʗ����_�w�}����Ӈ��@��U
��G��o�����W�W���������D�����g�b�o����9�ԜY�ƿ�T�������7�1�f�c�m��8���7���F��P ��U���&�2�7�1�d�h�MϜ�6����l�N�����u�%�&�2�5�9�D��CӤ��#��d��Uʦ�2�4�u�%�$�:����J���$��{+��N���u�&�2�4�w�-��������T�,��9���n�u�u�&�0�<�W���
����W��_��U�����n�u�w�.����Y����Z��S
��C���u����l�}�Wϭ�����R��^	�����c�u�u����L���Yӕ��]��V�����1�
�b�u�w��;���B�����Y�����<�
�1�
�o�}�W���5����9F������4�
�<�
�3��N���Y����v'��=d��Uʶ�8�:�0�!�:��@��@����U9��~=ךU���:�!�}�u�w�}�WϿ�&����	F��=��*����n�u�u�w�}����
����z(��c*��:���n�u�u�u�w�<�(�������z(��c*��:���n�u�u�u�w�<�(�������f2��c*��:���n�u�u�u�w�<�(�������f2��c*��:���n�u�u�u�w�<�(�������|3��d:��9����_�u�u�w�}��������l��T��;ʆ�������8���J�ƨ�D��^����u�u�u�;��3�������/��d:��9�������w�n�W������]ǻN��U���;��;�0�`�8�E��0�Ɵ�w9��p'��#����u�f�u�8�3���B���F���'���0�b�0�f�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����]9��Y	��B���a�o��u���8���&����|4�_�����:�e�n�u�w�}�WϷ�&����V9��R1�Oʜ�u��
����2���+������Y��E��u�u�u�u�>�����&Ĺ��F��~ ��!�����
����_������\F��d��U���u�<�
�4�0��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����4� �9�:�#�2�(������/��d:��9����_�u�u�w�}��������\��X��G���d�o��u���8���&����|4�_�����:�e�n�u�w�}�WϷ�&����R
��Y����
�
�u�u���3���>����F�N�����4� �9�:�#�2�(������/��d:��9�������w�n�W������]ǻN��U���;��;�4��3����H����F��~ ��!�����n�u�w�}�WϷ�&����R
��Y����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����R��[-�����
�g�0�c�m��W���&����p]ǻN��U���;��;�4��3����H����F��~ ��!�����
����_������\F��d��U���u�<�
�4�9��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����4�;�
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h)�����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����R��hZ��*���u������4���:����U��S�����|�_�u�u�w�}��������l��T��;ʆ�������8���J�ƨ�D��^����u�u�u�;��4�������/��d:��9�������w�n�W������]ǻN��U���;��<�&�c�8�A��0�Ɵ�w9��p'��#����u�f�u�8�3���B���F���2���&�a�0�b�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����]9��D��E���u��
���L���Y�����g8��*���u�u�����0���/����aF�N�����u�|�_�u�w�}�W���)����V9��N��U���
���
��	�%���Hӂ��]��G�U���u�u�<�
��o���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N�����
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƥ�l5��1��E���u��
���(���-��� W��X����n�u�u�u�w�4�(���H����\��yN��1��������}�D�������V�=N��U���u�%�'�!�%��W���,�Ɵ�w9��p'��#����u�f�u�8�3���B���F������'�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�W���YӇ��A��E ��U��� �u��
���(���-��� W��X����n�u�u�u�w�<�(�������\��b:��!�����
����_������\F��d��U���u�4�
�0�"�3�C��6����g"��x)��*�����}�d�3�*����P���F�N��*��� �;�`�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƭ�l��B��C��������4���:����U��S�����|�_�u�u�w�}��������F��x;��&���������W��Y����G	�UךU���u�u�%�'�#�/�(���Y����`2��{!��6�����u�f�w�2����I��ƹF�N�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����C9��T��;ʆ�����~�W�W����Ư�^��R ���ߊu�u�:�%�9�3�W���O����
 ��h��Dʜ�_�u�u�:�#�u�W���Y����C9��\N�<����
���l�}�W���YӇ��A��N��U���
���n�w�}�W�������R��N��U���
���n�w�}�W�������]�!��U���
���n�w�}�W�������_�!��U���
���n�w�}�W�������R��N��!ʆ�����]�}�W���Y����*��Y	��L���e�o��u���8���&����|4�_�����:�e�n�u�w�}�WϷ�&����R��hW��*���u������4���:����U��S�����|�_�u�u�w�}����
����\��yN��1�����_�u�w�}�W���)����Z��1��E���u��
���(���-��� W��X����n�u�u�u�w�4�(�������l^��h_��U���������4���Y����W	��C��\�ߊu�u�u�u�9������֓�lV�'��&���������W��Y����G	�UךU���u�u�;��>���������B9��T��;ʆ�������8���J�ƨ�D��^����u�u�u�;�3��W���7ӵ��l*��~-��0����}�d�1� �)�W���s���F�^ ����o��u����>���<����N��
�����e�n�u�u�w�}��������lV�!��U���
���
��	�%���Hӂ��]��G�U���u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�N�����0� �;�g�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���R��R����o������0���/����aF�N�����u�|�_�u�w�}�W�������z(��c*��:���u�n�u�u�2�9��������lǑN�����:�0�!�8��j�F���&ù��V��dd��Uʥ�'�u�_�u�w�}�W������/��d:��9����_�u�u�w�}��������}F��s1��2���_�u�u�u�w�-��������}F��s1��2���_�u�u�u�w�-����Y�ƃ�gF��s1��2���_�u�u�u�w�-����Y�ƃ�gF��s1��2���_�u�u�u�w�-���� ����f2��c*��:���n�u�u�u�w�4�(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����0� �;�e�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���R��R����o������0���/����aF�N�����u�|�_�u�w�}�W�������z(��c*��:���u�n�u�u�2�9��������lǑN�����:�0�!�8��j�F���&ù��W��B��G���f�;�
�g�d�;����
�ƅ�9F�	�����u�_�u�u�w�}�3��0����v4��N��U��������g�>���>����F�N�����
���u�w��2���B���F�
��D�����o����%�ԜY���F��B��<���u�u����}�L���YӖ��GF�N��U���6�>�o��w�	�(���0��ƹF�N�����u�u�����0���s���F�S��U���������!���6���F��@ ��U���_�u�u�u�w�4�F��0�Ɵ�w9��p'��#����u�f�u�8�3���B���F������o��u����>���<����N��S�����|�_�u�u�w�}���0�Ɵ�w9��p'�����u�u�u�:�#�g�8���*����|!��h8��!���}�d�1�"�#�}�^���s���V��T�����!�_�_�u�w�2�����ơ�rP��_��*ڊ�&�7�f�;��o���&����_
��D��&���u�2�;�'�4�u�W���Y����wF��~ ��2���_�u�u�u�w��(���>����z(��p+�����u�u�u�<�g�
�3���Cӯ��v!��d��U���u�1�;�
��	�W���7����a]ǻN��U���:�!����g�>���>���l�N�����_�u�u�u�w�1�W���7ӵ��l*��~-�U���u�u�'�&�#�g�>���-����t/��=N��U���u�<�e�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӂ��F��~ ��!�����
����_������\F��d��U���u�6�u�u���3���>����F�N�����u�u� �u���8���&����|4�_�����:�e�u�n�w�}��������]��dװU���6�8�:�0�#�0�6��H�ߪ�9��B��G���f�;�
�g�f�0����	ӯ��F�P�����}�u�u�u�w��W���7����a]ǻN��U��� �
���w�}�9���<��ƹF�N��������o��	�0���s���F�S��*����u�u����L���Y�����C1��1���o�����t�}���Y����NǻN��U���<�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������	F��=��*����
����u�FϺ�����O��N��U���1� �u�u��}�#���6����e#��x<��F���:�;�:�e�w�f�W�������\��Y��N�ߠ_�0�<�_�w�}����&ù�� 9��hX�U���:�%�;�;�w�m�A��Hʀ��l ��=N��U���!�8�%�}�w�}�W�������XF������_�u�u�u�w�-����D�ƭ�l��d��U���u�4�
�!�%�}�IϹ�	����l ��h��C���4�
�!�'�{�}�W���YӇ��W	��S����3�e�3�f�1��Fׁ�	����VJǻN��U���%�<�9�u�i�:����I����l ��_�����1�0�_�u�w�}�W�������[�P�����3�f�3�
�f���������F�N�����4�2�
�
��}�IϹ�	����l ��h��C���<�
�4�2���(��Y���F��Y1�����b�0�d�h�w�/�(���&����U��V�����;�0�b�0�f�W�W���Y�ƥ�l4��P��*���u�k�2�%�1�m��������9��h<�����
�
�y�u�w�}�WϷ�&����V9��R1�H���'�
�
�
�����A����a��R1����_�u�u�u�w�3�%����ѓ�lR�	N�����e�3�f�3��l�(���+����lQ��hZ�U���u�u�<�
�6�:�(؁�&�����h��*���
� �c�m�>�����&Ĺ��JǻN��U���;��;�0�`�8�A��Y����U9��Q1�����d�
�;��9�8�@���O���F�N��*���2�
�
�
�w�c�����֓�lU��B1�M���
�4�2�
���[���Y�����z�����;�'�9�d���W�������lV��h]�� ��m�<�
�4�"�1��������l��d��U���u�<�
�4�"�1��������l��S����3�e�3�f�1��Fׁ�����F��X �����g�0�d�_�w�}�W�������F��X �����g�0�g�h�w�/�(���&����U��V�����;�4��;�%�1�F݁�&��ƹF�N�����;�4��;�%�1�F݁�&�����h��*���
� �c�m�>���������A	��\��*���u�u�u�u�>���������A	��\��*���k�2�%�3�g�;�D���&����Z��V �����!�:�
�g�2�i�}���Y���Z��V �����!�:�
�g�2�h�J�������9��1��*��
�;��;�6���������V9��=N��U���u�;��;�6���������V9��
P�����
�
�
�
�"�k�O���&����R
��Y����
�
�y�u�w�}�WϷ�&����R
��Y����
�
�u�k�0�-�����Փ�F9��1��*��� �9�:�!�8��E���N���F�N��*���;�
�
�
�w�c�����֓�lU��B1�M���
�4�;�
���[���Y�����p�����0�d�h�u�%��(߁�&����lP��h��2���&�a�0�d�]�}�W���Y����R��hZ��*���k�2�%�3�g�;�D���&����Z��V��*ފ�
�y�u�u�w�}��������9��N��U���
�
�
�
��(�A�������Z��1��F�ߊu�u�u�u�9�����M����[�P�����3�f�3�
�f���������l��d��U���u�<�
�4�9��(���Y����A��h^��*ي� �c�m�<��<����&����9F�N��U����<�&�a�2�k�J�������9��1��*��
�;��<�$�i���s���F�^ �����
�
�
�u�i�:����I����l ��_�����4�;�
�
��q�W���Y����]9��D��E��u�'�
�
���(���O�ޓ�]9��D��E�ߊu�u�u�u�9��(݁�&�����h��*���
� �c�m�>��!�������F�N������g�0�d�j�}����&ù�� 9��hX�*����
�
�
�{�}�W���Yӏ��c0��h��U��2�%�3�e�1�n����H˹��l6��1��G�ߊu�u�u�u�9��(݁�&�����h��*���
� �c�m�>��!�������F�N������d�0�e�j�}����&ù�� 9��hX�*����
�
�
�{�}�W���Yӏ��`6��h��U��2�%�3�e�1�n����H˹��l5��1��D�ߊu�u�u�u�'�/����&�����h��*���
� �c�m�6���������F�N�����0� �;�d�j�}����&ù�� 9��hX�*���'�!�'�
�{�}�W���YӇ��A��E ��U��2�%�3�e�1�n����H˹��l��B��G�ߊu�u�u�u�'�/����&�����h��*���
� �c�m�6���������F�N�����0� �;�a�j�}����&ù�� 9��hX�*���'�!�'�
�{�}�W���YӇ��A��E ��U��2�%�3�e�1�n����H˹��l��B��@�ߊu�u�u�u�'�/����&�����h��*���
� �c�m�6���������F�N�����0� �;�b�j�}����&ù�� 9��hX�*���'�!�'�
�{�}�W���YӇ��A��E ��U��2�%�3�e�1�n����H˹��l��B��M�ߊu�u�u�u�'�/����&�����h��*���
� �c�m�6���������F�N�����0�h�u�'���(���&����^��G1��\�ߠu�u�2�%�1�m���&����W������;�u�e�c�b�l��������F�G��U���u�_�u�u�w�}�������R��[�U���u�u�4�
�$�}�IϿ�&����9F�N��U���&�4�!�h�w�/�(���&����l ��X�����!�'�y�u�w�}�WϿ�&����[�P�����3�d�
� �a�l��������F�N�����1�0�h�u�%��(߁�&�ד�F9��1��*���0�_�u�u�w�}�������F��G1��E���d�
� �c�f�<�(�����ƹF�N������4�2�
���W�������lV��h_�����c�
�;���<����&����9F�N��U�����4�2���(���GӁ��l ��h��D���
�c�
�;������&ʹ��JǻN��U���;�'�&�!�c�`�W���&����U9��h��C���<�
�0�0��q�W���Y����]9��{	�����
�
�u�k�0�-��������U��_������4�;�
���[���Y�����g"�����
�
�
�u�i�:����I����9��hX�*�����4�;���(��Y���F��Y1�����;�e�0�e�j�}����&ù��W��B1�D���
�!�!����(��Y���F��Y1�����%�6�0��2��B��Y����U9��Q1�*���c�d�<�
�%�9��������V��BךU���u�u�;�1��}�IϹ�	����l ��1��*��
�;�1�
�{�}�W���Yӏ��e��S����3�e�3�d��(�A�������lU�N��U���4�
�0� �9�m�J�������9��_�� ��d�4�
�0�"�3�G�ԜY���F��h�� ���d�h�u�'���(���H����P��V�����;�d�_�u�w�}�W�������]9��
P�����
�
�
�d�1��Aށ�	����F��BךU���u�u�%�'�#�/�(���GӁ��l ��h��D���
�c�
�%�%�)����U���F������k�2�%�3�g�;�Fށ�����l��T����u�2�%�3�g�;�F߁�����\��X�����u�e�c�`�f�;�G���H���F��E�����_�u�u�u�w�-����D�ƭ�l��d��U���u�4�
�&�w�c����
��ƹF�N�����4�!�h�u�%��(߁�&�֓�F9��1��*���'�y�u�u�w�}�������F��G1��E���d�
� �c�o�<�(������F�N��*���0�h�u�'���(���I����Q��V�����_�u�u�u�w�-���� ���T��Q1����
� �c�m�6�����U���F�����h�u�'�
���(�������9��h��Y���u�u�u�4��8����I���T��Q1����
� �c�m�6���������F�N�����0� �;�d�j�}����&ù��V��B1�M���
�0� �;�f�W�W���Y�ƭ�l��
P�����
�
�
�e�1��@ׁ�	����lǻN��*ڊ�4�1�&�7�d�3�(���
���� 9��[�����c�u�u�:�'�3����I����W��h^�����&�7�f�;��o���&����_
��DךU���0�0�<�u�6�}�}���Y���z"�	N����u�u�u� ��	�0���G����F�N�����
���u�i�n�[���Y�����1��1���h�u�g�_�w�}�W�������z"��S�F���u�u�%�'�w�<�W�ԜY���F��\N��U���6�>�_�u�w�}�W��������E�����u�u�u�<�g�`�W���&����Q��BךU���u�u�<�d�j�}��������l��=N��U���u�%�:�0�j�}��������l	��X
�����u�u�u�0�j�}��������l��=N��U���u�:�!�h�w�/�(���O�ѓ�O��=N��U���
�4�1�&�5�n����K����9��Q��*���
�c�u�u�8�-����Y�֍�S����*���1�&�7�f�9��E���J����U��h
�����u�0�0�<�w�<�W�ԜY���F��S�D�ߊu�u�u�u���#���Y���l�N��Uʱ�;�
���w�c�D��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��|�u�u�%�%�}����s���F�T��H���%�6�>�_�w�}�W�������X��G1���ߊu�u�u�u�>�m�J�������lP��h����u�u�u�<�f�`�W���&����
W��BךU���u�u�%�:�2�`�W���&����
W��G���ߊu�u�u�u�2�`�W���&����
W��RBךU���u�u�:�!�j�}��������l��dךU���
�
�&�7�d�3�(���
���� 9��[�����c�u�u�:�'�3����I����W��h^�����f�;�
�g�$�n�(܁�����@ǻN�����<�u�4�u�]�}�W���Y���F��=N��U���u� �
���}�I��s���F�S��*����u�k�f�{�}�W���Yӂ��9��s:��H���g�_�u�u�w�}����.����[�\��U���%�'�u�4�w�W�W���Y�Ư�XF������_�u�u�u�w�8����GӇ��A��=N��U���u�<�e�h�w�/�(���O�ӓ�JǻN��U���<�d�h�u�%����L����9F�N��U���h�u�'�
�"�k�B���U���F�
����u�'�
� �a�h����s��� ��h����;�
�g�&�d��(�������l3��T�����;�;�u�e�a�h�Fָ�I����Q9��Y��G���f�
�
� �;�9����YӁ��V����U�ߊu�u�u�u��`�W��Y���F��b#��!���u�k�f�_�w�}�W����֓�z"��S�F���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���K���F��E�����_�u�u�u�w�1�W�������XJǻN��U���0�0�u�k�6����Y���F��^ �H���'�
� �c�n�-�[���Y�����N��U���
� �c�l�'�q�W���Y����VF�	��*���c�l�6�y�w�}�W�������X��E�� ��l�%�|�_�w�}�������� T��h]����
�
�4�
�$��A���Y����\��CN��4��d�l�
�
�:�1�Dݰ�&�Ԣ�lU��1�����%�u�u�2�9�/�ϳ�	��ƹF�N��1��u�y�u�u�w�}�9���*����[�BךU���u�u�<�e� ��?��Y����F�N�����
���u�i�n�[���Y�����C1��1���h�u�g�_�w�}�������9F�N��U���e�h�u�'��(�@���	��ƹF�N����h�u�'�
�"�j�@���U���F�
����u�'�
� �`�j����s��� ��h����;�
�g�&�d��(���&����fP��N�����0�!�8��`�l�N���&����lU��D1����g�d�8�-�3�-�W�������Z��V�����u�u�u��j�}�[���Y���(��h=��2���k�d�_�u�w�}�W���I����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���:�!����`�W��s���C	����U�ߊu�u�u�u�>�m�J�������lQ��h����u�u�u�<�f�`�W���&����T��BךU���u�u�:�!�j�}��������l��dךU���
�
�8�9�d�3�(���
����9��O1�����b�o�6�8�8�8�ϳ�8����_��1�� ���g�&�f�;��o�F�������9F�	�����u�4�u�_�w�}�W���=���JǻN��U��� �
���w�c�F�ԜY���F��Y^��<���u�k�f�y�w�}�W�������d/��N��U��_�u�u�u�w�2����=���F��d��Uʥ�'�u�4�u�]�}�W���Y����[�P�����d�
�e�_�w�}�W������F��G1��*��
�d�_�u�w�}�W������T��Q��D݊�g�n�_�u�w��(�������@9��Y��G���8�-�1�%��e�MϽ�����]��/�@��3�e�3� ��o�������lW��V���ߊu�u�0�0�>�}����s���F�~*��K��_�u�u�u�w��(���>���W�N��U���1�;�
���}�I��U���F�
��D�����h�u�e�W�W���Y�ƨ�F��~*��U��f�|�u�u�'�/�W���Y���F�N�����k�2�%�3��o�(��s���F�S��U��2�%�3�
�e��F�ԜY���F��B��Kʲ�%�3�
�g��o�L�Զs���F���U���'�;�u�!�#�}����*����F����U���!�u�4�=�9�s�Z�ԜY�ƭ�l%��Q�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�u�u�w�}�W���Y���F���6���&�u�h�4������s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�'���(���I����Q��V�����
�%�&�4�#�/�Ͽ�
����C��R��U���u�u�2�%�1�m���&����^��G1�����4�
�!�'��8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���T��Q1����
� �c�m�6�����&����G��h��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9�� 1����|�u�=�;�]�}�W���Y���F�N�����3�e�3�d��(�A�������R��V�����
�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�1����Q����\��h�����u�u�'�
���(�������9��h�����u�=�;�_�w�}�W���Y���F�N�����e�3�d�
�"�k�O���&����G9��h�����0�u�h�4��2��������]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����֓�lW��Q��Cۊ�%�&�4�!�6�����&����R��P �����&�{�x�_�w�}����&ù��W��B1�D���
�!�'�
�'�.��������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N�����
�
�
�d�1��Aށ�	����A��G1�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���f�3�8�d�~�t����Y���F�N��U���u�u�u�'���(���H����P��V�����
�%�&�4�#�/���Y����\��h�����n�u�u�u�w�}�W���YӃ��Z ������!�9�2�6�f�`�����֓�lW��Q��Cۊ�%�'�4�,�~�)����Y���F�N��U���u�u�'�
���(�������9��h�����%�&�4�!�%�:�K���	����@��X	��*��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���T��Q1�����3�
�d�
�'�.��������R��E�����2�u�'�6�$�s�Z�ԜY�ƫ�C9��1��F���
�d�
�%�$�<����&����G9��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�2�%�3�g�;�D���&����R��C��*���&�4�!�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�a�1�0�F�������\�V�����
�:�<�
�w�}����&ù��W��B1�D���
�:�0�|�~�)����Y���F�N��U���u�u�'�
���(܁�����l��D�����
�!�'�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�w�}�W�������N��h�����:�<�
�u�w�/�(���&����U��V�����4�,�|�!�2�}�W���Y���F�N��U���'�
�
�
�����A����@��C1��*���'�
�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	����`��X�����e�4�
�9��/�Ͽ�
����C��R��U���u�u�%�d��8��������9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�F߁�����]��R1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��G���8�g�|�u�?�3�}���Y���F�N��U���u�u�%�d��8��������9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��E���!�0�u�u�w�}�W���Y���F�N��U���e��!�:�9�.��������W9��R	��Hʥ�d�
�0�%�>�)�(���&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�l�(���	����@9��1�����&�<�;�%�8�8����T�����1�����;�&�0�e�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��h=�����!�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�Hù��G��Y�����4�
�9�|�~�)����Y���F�N��U���u�u�
�e��)����
����l��PN�U���e��!�:�9�.���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
�f�����&����R��[
�����4�&�2�u�%�>���T���F��_�����&�0�e�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���D���%�!�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����H����[��=N��U���u�u�u�u�w�}�W���Y����l/��B�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�g�~�)����Y���F�N��U���u�u�u�u��l�>�������9��h��*���2�i�u�
�f�����&����R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p���&����G��h^�����4�&�2�u�%�>���T���F��_�����&�0�e�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�W��Y�����e�%�0�u�j�<�(���
���� T��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��F���	����V9��V�����|�!�0�u�w�}�W���Y���F�N��*����%�!�
������E�Ƽ�W��Y�����e�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h_��<���!�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��F���	����V9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}���&����G��h_�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�d�|�!�2�}�W���Y���F�N��U���u�u�
�d��-����&¹��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��\�����u�u�u�u�w�}�W���Y���F���D���%�!�
�
��-����	����[��h_��<���!�
�
�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�d�
�;� �$�8�F����ƭ�@�������{�x�_�u�w��F���	����V9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
�f�����&����C��R�����:�&�
�#�e�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*����%�!�
���������G��d��U���u�u�u�u�w�}�WϮ�H¹��C��h��*���2�i�u�
�f�����&����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�Fށ�����l��h�����%�0�u�&�>�3�������KǻN��*����%�!�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�d�
�;� �$�8�E���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����1�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�i�F������F�N��U���u�u�u�u�w�}���&����G��h\�����1�%�0�u�j�-�Fށ�����l��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����l/��B�����%�0�u�&�>�3�������KǻN��*����%�!�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h_��<���!�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�H¹��C��h��*���#�1�|�u�?�3�}���Y���F�N��U���%�d�
�;�"�.����	����[��h_��<���!�
�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C���
�;� �&�2�n��������V��D��ʥ�:�0�&�u�z�}�WϮ�H¹��C��h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����l/��B�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���g�3�8�g�~�}����s���F�N��U���u�u�u�u�'�l�(�������lU��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��A��u�=�;�_�w�}�W���Y���F�N��Uʥ�d�
�;� �$�8�D���&����C��R����
�;� �&�2�n������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�d��-����&����V��D��ʥ�:�0�&�u�z�}�WϮ�H¹��C��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�Fށ�����l��h����u�%�6�;�#�1�D݁�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�d�
�;�"�.��������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�W��Y�����f�%�0�u�j�-�Fށ�����l��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&�ד�]��D1��A���
�9�
�'�0�<����Y����V��C�U���%�d�
�;�"�.��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�d��-����&ǹ��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��_��U���;�_�u�u�w�}�W���Y���F�N��Dۊ�;� �&�0�c�<�(���&����Z�V�����
�:�<�
�l�}�W���Y���F�N��U���<�u�4�
�>�����L����[��=N��U���u�u�u�u�w�}�W���Y����l/��B�����4�
�9�
�%�:�K���&�ד�]��D1��A���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����1�����
�
�
�'�0�<����Y����V��C�U���%�d�
�;�"�.����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N����
�;� �&�2�i����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�W��Y�����a�4�
�9�~�t����Y���F�N��U���u�u�u�
�f�����&����C��R����
�;� �&�2�i�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�d��'�)�(���&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�W��Y�����`�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����1�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��F�������9F�N��U���u�u�u�u�w�}�W���H����F��R1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�c�|�!�2�}�W���Y���F�N��U���u�u�
�d��-����&ƹ��l��h����u�
�d��'�)�(���&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�l�(�������lS��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�W��Y�����`�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&�ד�]��D1��@���0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
�f�����&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h_��<���!�
�
�
�%�:�K���&�ד�]��D1��@�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lW��~ �����
�
�%�#�3�-����
������T��[���_�u�u�
�f�����&����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�l�(�������lP��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�d��%�#��(ف�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������Q�C��U���u�u�u�u�w�}�W���Y�����1�����
�
�
�%�!�9����Y����lW��~ �����
�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��Dۊ�;� �&�0�a�-����
������T��[���_�u�u�
�f�����&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�d��'�)�(���&����Z�V�����
�#�g�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h_��<���!�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�Fށ�����l��h����u�
�d��'�)�(���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�c�����:����\
��h^�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�4� �9�8�)����&ù��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�c�����:����\
��h^�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�d�|�!�2�}�W���Y���F�N��U���u�u�
�
�6�(��������V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��u�=�;�_�w�}�W���Y���F�N��Uʥ�a��;�4��3�����֓�C9��S1�����h�%�a��9�<�4�������lV��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ǹ��]��t�����0�e�%�0�w�.����	����@�CךU���
�
�4� �;�2����&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�4�"�1��������9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�%�c�����:����\
��h^�����1�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G��U���;�_�u�u�w�}�W���Y���F��1������;�'�9�2�m����Y����lR��V �����!�:�
�
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�a��;�4��3�����ד�C9��S1�����&�<�;�%�8�8����T�����h#�� ���:�!�:�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�a��;�4��3�����ד�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h\�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ފ�4� �9�:�#�2�(���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lW��N�����u�u�u�u�w�}�W���Y���F��hZ�����9�:�!�:���(�������A��S��*ފ�4� �9�:�#�2�(���&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�i�:�������G��h��*���2�4�&�2�w�/����W���F�G1��8���4��;�'�;�8�F�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��A���;�4��;�%�1����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1������;�'�9�2�l���������YNךU���u�u�u�u�w�}�W���&ǹ��]��t�����0�d�%�0�w�`����4����_%��C��*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1������;�'�9�2�o��������V��D��ʥ�:�0�&�u�z�}�WϮ�M����F��X �����
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1������;�'�9�2�o��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�E�������F��R ��U���u�u�u�u�w�}�W���Y����lR��V �����!�:�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���O�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ғ�R��[-�����
�
�
�%�!�9����Y����lR��V �����!�:�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�a��;�6���������l��PN�����u�'�6�&�y�p�}���Y����~��V�����9�0�g�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��Y��6���'�9�0�g�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ғ�R��[-�����
�
�
�%�!�9�^������F�N��U���u�u�u�u�'�i�:�������G��h��*���2�i�u�
��<��������_9��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ғ�R��[-�����
�
�
�%�!�9����Y����T��E�����x�_�u�u����������A	��R1�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ғ�R��[-�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��F�������9F�N��U���u�u�u�u�w�}�W���&����R
��Y�����f�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�e�t����Y���F�N��U���u�u�u�u�w��(�������]��[1��F���
�9�
�'�0�a�W���&����R
��Y�����f�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*��� �9�:�!�8��(܁�����@��YN�����&�u�x�u�w�-�C�������\��X��*ي�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����4����_%��C��*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�i�:�������G��h��*���#�1�|�u�?�3�}���Y���F�N��U���%�a��;�6���������l��PN�U���
�4� �9�8�)����&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�i�:�������G��h��*���#�1�%�0�w�.����	����@�CךU���
�
�4� �;�2����&����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�i�:�������G��h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��G؊�&�
�d�|�#�8�W���Y���F�N��U���u�u�u�
��<��������_9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����f�|�!�0�w�}�W���Y���F�N��U���u�
�
�4�"�1��������9��h��*���2�i�u�
��<��������_9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l+��B�����:�
�
�
�%�:�����Ƽ�\��D@��X���u�%�a��9�<�4�������lR��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�a��3��������l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�4�"�1��������9��h��\���!�0�u�u�w�}�W���Y���F���*��� �9�:�!�8��(ہ����F��1������;�'�9�2�i�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�4�"�1��������9��h��*���2�4�&�2�w�/����W���F�G1��8���4��;�'�;�8�B���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�4�"�1��������9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���u�=�;�_�w�}�W���Y���F�N��Uʥ�a��;�4��3�����ӓ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��Z�U���;�_�u�u�w�}�W���Y���F�N��A���;�4��;�%�1��������W9��R	��Hʥ�a��;�4��3�����ӓ�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ہ�����p	��E�����%�0�u�&�>�3�������KǻN��*ފ�4� �9�:�#�2�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�4� �9�8�)����&ƹ��V�
N��*���&�
�#�g�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*��� �9�:�!�8��(ځ�	����O�C��U���u�u�u�u�w�}�W���YӖ��l+��B�����:�
�
�
�%�:�K���&ǹ��]��t�����0�`�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*��� �9�:�!�8��(ف�	����l��PN�����u�'�6�&�y�p�}���Y����~��V�����9�0�c�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*��� �9�:�!�8��(ف�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����W����ߊu�u�u�u�w�}�W���Y���F��1������;�'�9�2�k��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��Y��6���'�9�0�c�6��������F��1������;�'�9�2�k������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�(��������V9��G��U���<�;�%�:�2�.�W��Y����lR��V �����!�:�
�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h#�� ���:�!�:�
������E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��Y��6���'�9�0�c�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(ہ�����p	��E�����%�0�u�h�'�i�:�������G��h��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Y��6���'�9�0�b�6���������@��YN�����&�u�x�u�w�-�C�������\��X��*݊�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��Y��6���'�9�0�b�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!�e�;���P�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ғ�R��[-�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�l�F������F�N��U���u�u�u�u�w�}����4����_%��C��*���
�%�#�1�'�8�W��	�ғ�R��[-�����
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����;�4��9�/����N����TF��D��U���6�&�{�x�]�}�W���&����R
��Y�����b�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ǹ��]��t�����0�b�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ہ�����p	��E�����4�
�9�|�~�)����Y���F�N��U���u�u�
�
�6�(��������V9��G��U��%�a��;�6���������l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ځ�����V9��V�����'�2�4�&�0�}����
���l�N��@���;�0�0�e�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�4�2�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����H����[��=N��U���u�u�u�u�w�}�W���Y����a��R1��E���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�}�W���YӃ��Z �V�����1�
�b�|�#�8�W���Y���F�N��U���u�u�u�
��<����&ù��l��h����u�
�
�4�0��(߁�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�b������֓�A��V�����'�6�&�{�z�W�W���&ƹ��]��R1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������9��R	��Hʴ�
�:�&�
�!�o�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�4�2�
���������G��d��U���u�u�u�u�w�}�WϮ�L����T��h^�����i�u�
�
�6�:�(���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�b������ד�C9��S1�����&�<�;�%�8�8����T�����h<�����
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����0�d�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�o�^������F�N��U���u�u�u�u�w�}����+����l��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����l�u�=�;�]�}�W���Y���F�N��U���%�`��;�2�8�F���&����C��R������;�0�0�f�<�(���B���F�N��U���u�u�u�;�w�;�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�4�0��(ށ�����@��YN�����&�u�x�u�w�-�B�������lW��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�`��3����H����TF������!�9�f�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��'���0�0�d�4��1�^�������9F�N��U���u�u�u�u�w��(�������9��R	��Hʥ�`��;�0�2�l�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�4�0��(݁�	����l��PN�����u�'�6�&�y�p�}���Y����a��R1��G���
�9�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l4��P��*؊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�)����Y���F�N��U���u�u�u�u������&����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��h_�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ߊ�4�2�
�
��-����	����[��h[�����
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����;�0�0�e�-����
������T��[���_�u�u�
��<����&����V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�4�2���(������R��X ��*���g�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lS��V ��*���
�%�#�1�~�}����s���F�N��U���u�u�%�`��3����K����TF���*���2�
�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����;�0�0�d�<�(���&������^	�����0�&�u�x�w�}����+����l��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����V9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C\�����g�|�u�=�9�W�W���Y���F�N��U���u�%�`��9�8��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����_�����ߊu�u�u�u�w�}�W���Y���F��1�����0�f�4�
�;�����E�Ƽ�9��Y	�����4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h[�����
�
�
�'�0�<����Y����V��C�U���%�`��;�2�8�D�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��@���;�0�0�f�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ƹ��]��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�4�2���(������C9��e�����f�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h[�����
�
�
�%�!�9����Y����T��E�����x�_�u�u������&����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�h�%�������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���!�0�u�u�w�}�W���Y���F�N��U���
�4�2�
����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����K���G��d��U���u�u�u�u�w�}�W���YӖ��l4��P��*ފ�%�#�1�%�2�}�JϮ�L����T��hZ�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Y	�����%�0�u�&�>�3�������KǻN��*ߊ�4�2�
�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h<�����
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�B�������lR��G1�����u�=�;�_�w�}�W���Y���F�N��@���;�0�0�a�'�8�W��	�ӓ�R��h��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Y	�����4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�`��9�8��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�6�:�(���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���K����^9��G�����_�u�u�u�w�}�W���Y���F�G1��'���0�0�`�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��F�������9F�N��U���u�u�u�u�w�}�W���&����V9��1��*���
�'�2�i�w��(�������9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L����T��h[�����4�&�2�u�%�>���T���F��1�����0�`�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����a��R1��@���0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��<����&ƹ��l��G�����u�u�u�u�w�}�W���Y�����h<�����
�
�'�2�k�}�(ځ�����V9��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L����T��hX�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�4�2�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�`��;�0�2�k��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�E�������F��R ��U���u�u�u�u�w�}�W���Y����lS��V ��*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�g�c�}����s���F�N��U���u�u�u�u�'�h�%�������l��A�����u�h�%�`��3����O����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(�������9��R	�����;�%�:�0�$�}�Z���YӖ��l4��P��*܊�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����+����l��h����u�%�6�;�#�1�D݁�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�`��;�2�8�A���&����O��_�����u�u�u�u�w�}�W���Y����a��R1��C���0�u�h�%�b���������F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(�������9��h��*���2�4�&�2�w�/����W���F�G1��'���0�0�b�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���2�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�g��.�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ƹ��]��R1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
�6�:�(���&����_��E��I���
�
�4�2���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`��3����N����TF��D��U���6�&�{�x�]�}�W���&����V9�� 1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u������&����C��R�����:�&�
�#�e�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ߊ�4�2�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����+����l��h����u�
�
�4�0��(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`��3����A����E
��G��U���<�;�%�:�2�.�W��Y����lS��V ��*���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��e�����m�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�e�t�W������F�N��U���u�u�u�u�w�-�B�������l^��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��G��u�=�;�_�w�}�W���Y���F�N��Uʥ�`��;�0�2�e��������V�
N��@���;�0�0�m�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�4�2���(���Ӈ��Z��G�����u�x�u�u�'�h�%�������l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�`��9�8����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����0�m�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u������&����C��R������;�0�0�o�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�4�2���(�������A��V�����'�6�&�{�z�W�W���&ƹ��]��R1�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ӓ�R��h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��G؊�&�
�d�|�#�8�W���Y���F�N��U���u�u�u�
��<����&ʹ��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��_�����u�u�u�u�w�}�W���Y���F���*���2�
�
�
�'�+���������h<�����
�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��@���;�0�0�l�'�8�W�������A	��D�X�ߊu�u�
�
�6�:�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�4�2�
������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l4��P��*ӊ�%�#�1�|�w�5��ԜY���F�N��U���u�%�`��9�8����	����[��h[�����
�
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��C���'�8�!�'���(�������A��V�����'�6�&�{�z�W�W���&Ź��A��C��*���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��g�����'�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�g��.�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ź��A��C��*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�g�g�}����s���F�N��U���u�u�u�u�'�k�'�������@9��1��*���
�'�2�i�w��(�������A��h^�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��E�����
�
�
�'�0�<����Y����V��C�U���%�c��'�:�)����&ù��V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�4�4�2�8����I����TF������!�9�f�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��%���8�!�'�
���������G��d��U���u�u�u�u�w�}�WϮ�O����R��R�����%�0�u�h�'�k�'�������@9��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�Г�R��R�����d�4�
�9��/�Ͽ�
����C��R��U���u�u�%�c��/��������9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�A�������V��R1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��G���8�g�|�u�?�3�}���Y���F�N��U���u�u�%�c��/��������9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��C���!�0�u�u�w�}�W���Y���F�N��U���
�4�4�0�2�.��������W9��R	��Hʥ�c��'�8�#�/�(���&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�k�'�������@9��1�����&�<�;�%�8�8����T�����h>�����0�&�0�d�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��g�����'�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�O����R��R�����4�
�9�|�~�)����Y���F�N��U���u�u�
�
�6�<����
����l��PN�U���
�4�4�0�2�.���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��<����&ù��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��p�����e�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h)�����
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�4�;���(�������A��S��*݊�4�;�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b��<�$�8�G����ƭ�@�������{�x�_�u�w��(�������9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�6�3�(���&����Z�V�����
�#�g�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY�����
�
�
�%�!�9�^������F�N��U���u�u�u�u�'�j�0���
����l��PN�U���
�4�;�
��f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b��<�$�8�F���&����C�������%�:�0�&�w�p�W���	�ѓ�R��h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����t��D1��D���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�w�5��ԜY���F�N��U���u�u�u�%�`������ד�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��^�U���;�_�u�u�w�}�W���Y���F�N��B���<�&�0�d�6��������F�� 1�����0�d�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��/�Ͽ�
����C��R��U���u�u�%�b��4����H����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��<�&�2�l����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��^ �����4�
�9�|�~�)����Y���F�N��U���u�u�
�
�6�3�(���&����Z�G1��2���&�0�d�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-����	����R��P �����&�{�x�_�w�}�(؁�����V9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����>����l��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y�����T�����2�6�d�h�6�����
����g9��\�����d�|�!�0�w�}�W���Y���F�N��U���u�
�
�4�9��(݁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������S�C��U���u�u�u�u�w�}�W���Y�����h)�����
�
�%�#�3�-����DӖ��l!��Y��*؊�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�����0�g�%�0�w�.����	����@�CךU���
�
�4�;���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���;�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N����]��h\�����1�|�u�=�9�W�W���Y���F�N��Uʥ�b��<�&�2�o����Y����lQ��V��*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�����0�f�4�
�;���������]F��X�����x�u�u�%�`������Փ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u������&����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���F�N������<�&�0�d�<�(���&����Z�V�����
�:�<�
�l�}�W���Y���F�N��U���<�u�4�
�>�����K����[��=N��U���u�u�u�u�w�}�W���Y����t��D1��F���
�9�
�'�0�a�W���&����@9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ي�'�2�4�&�0�}����
���l�N��B���<�&�0�f�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��p�����f�%�0�u�j�<�(���
���� T��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(������� 9��h��\���!�0�u�u�w�}�W���Y���F���*���;�
�
�
�%�:�K���&Ĺ��Z��R1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ފ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�4�9��(ہ�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�b��>�.��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���K����lT��N�����u�u�u�u�w�}�W���Y���F��hY�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�n�D������F�N��U���u�u�u�u�w�}����>����l��h�����%�0�u�h�'�j�0���
����l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����@9��1�����&�<�;�%�8�8����T�����h)�����
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ѓ�R��h��*���2�i�u�%�4�3����J����9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�b��4����M����E
��G�����_�u�u�u�w�}�W���Y���C9��p�����a�%�0�u�j�-�@�������lR��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����@9��1��*���
�'�2�4�$�:�W�������K��N������<�&�0�b�<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�4�;�
����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�}�'�>��������lW������6�0�
��$�o�(���&�����YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��^ �����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�a�~�)����Y���F�N��U���u�u�u�u������&����R��[
�����i�u�
�
�6�3�(���&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�j�0���
����l��PN�����u�'�6�&�y�p�}���Y����t��D1��@���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�4�;���(������F��R ��U���u�u�u�u�w�}�W���	�ѓ�R��h��*���2�i�u�
��<����&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�j�0���
����l��A�����u�&�<�;�'�2����Y��ƹF��hY�����
�
�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��2���&�0�c�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�g�1�0�E���Y����l�N��U���u�u�u�u�w�}�WϮ�N����]��hX�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����f�d�u�=�9�W�W���Y���F�N��U���u�%�b��>�.��������W9��R	��Hʥ�b��<�&�2�k������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�3�(���&������^	�����0�&�u�x�w�}����>����l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`������Г�A��S�����;�!�9�f��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��B���<�&�0�c�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(؁�����V9��G��U��%�b��<�$�8�A�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�3�(���&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��V��*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�f�t����Y���F�N��U���u�u�u�u�w��(�������9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��C���!�0�u�u�w�}�W���Y���F�N��U���
�4�;�
����������TF���*���;�
�
�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�b��<�&�2�j����Y����T��E�����x�_�u�u������&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�4�9��(؁����F��h�����#�g�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h)�����
�
�%�#�3�t�W������F�N��U���u�u�u�%�`������ѓ�A��S��*݊�4�;�
�
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�b��<�&�2�e��������V��D��ʥ�:�0�&�u�z�}�WϮ�N����]��hV�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��Z��R1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��G���8�g�|�u�?�3�}���Y���F�N��U���u�u�%�b��4����A����E
��G��U��4�
�:�&��2����B���F�N��U���u�u�u�9�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��2���&�0�m�4��1�(������C9��p�����m�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���;�
�
�
�%�:�����Ƽ�\��D@��X���u�%�b��>�.����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������<�&�0�o�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����t��D1��M���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�4�9��(ׁ����F�� 1�����0�m�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���;�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(�������
9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�@�������l_��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�4�;���(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lQ��V��*���
�%�#�1�'�8�W��	�ѓ�R��h��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��p�����l�%�0�u�$�4�Ϯ�����F�=N��U���
�4�;�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hY�����
�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����>����l��h�����|�u�=�;�]�}�W���Y���F�N������<�&�0�n�-����DӖ��l!��Y��*��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��d�����0�e�4�
�;���������]F��X�����x�u�u�%�n�����
����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�l��2�6�.��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&���� ^�����ߊu�u�u�u�w�}�W���Y���F��1�����&�0�e�4��1�(������C9��d�����0�e�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ӊ�<�;�9�
����������]F��X�����x�u�u�%�n�����
����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�l��0�<����I����TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���;�9�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����*����_��h^�����i�u�
�
�>�3����&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�d�$�������lW��G1�����0�u�&�<�9�-����
���9F���*���;�9�
�
��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������2�4�&�2�l��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�E�������F��R ��U���u�u�u�u�w�}�W���Y����l_��^	�����
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W���Y���F��D��]���&�2�7�1�d�k�W������F�N��U���u�u�u�u�w�-�N�������l��h�����%�0�u�h�'�d�$�������lW��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ʹ��T��D1��D���0�u�&�<�9�-����
���9F���*���;�9�
�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h=�����
�
�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R
��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�<�;�;��(ށ����F��1�����&�0�d�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����;�%�:�0�$�}�Z���YӖ��P��F��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y�����Yd��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���������� O��Y
�����4�
�:�&��2����Y�ƫ�C9��1��Dۊ� �c�d�4��2����PӒ��]l�N��U���u�u�u�6���3���2����F�� 1����i�u�'�
���(�������9��h�� ���e�_�u�u�w�}�W���Y�Ư�l��R1�����=�0��4�2��(���&¹��T9��^��Hʲ�%�3�e�3�f����H����A��E ��N���u�u�u�u�w�}�WϽ�&����l��Z1�����=�&���$�>�E�������F�	��*���
�
�d�3��k�(�������]9��=N��U���u�u�u�u�w�����&����l2��R������
�'�
�2��@��E�ƫ�C9��1��Dۊ� �c�d�4��8����J���F�N��U���u�3�
������&¹��T9��V��Hʲ�%�3�
�m��o�}���Y���F�N��������!��?����&�ޓ�l��h_�A��u�'�
� �a�l���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��B���8�c�|�u�?�3�W���Y���F�N��������:�#�(�(����֓�V��Z�I���9�����2����&�ѓ�l��d��U���u�u�u�u�w�;�(���;����lW��1����`�u�h�2�'�;�(��&����F�N��U���u�u�3�
���8���K����A��X�U��2�%�3�
�n��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��@���8�d�|�4�3�3����	����@��X	��*���u�'�
�
���(���O�ޓ�C9��Y��\���=�;�u�u�w�}�W���Y����_9��S������&�4�0��3����
�ד�V�� \�I���'�
�
�
�����A����A��E ��N���u�u�u�u�w�}�WϽ�&����l��Z1�����0��;�'�;�.�E�������F�	��*���
�
�
� �a�e��������lT��N��U���u�u�u�u�4���������p��V
��6���'�9�&�f�%�:�F��Y����A��h^��*ي� �c�m�4��8����J���F�N��U���u�6�
�:�2�)��������V��Y�����a�'�2�d�d�}�JϹ�	����l ��h��C���4�
�0� �9�i�}���Y���F�N�����:�0�!�'��<��������A	��D1�����d�a�u�h�0�-�����Փ�F9��1��*��� �;�`�_�w�}�W���Y���F��h �����'�
�4�6�3�9��������9��P1�A���h�2�%�3�g�;�D���&����R��R����_�u�u�u�w�}�W���Y����\��C��*���6�1�1�:�#�2�(���&����Q��R�����3�e�3�f�1��Fׁ�	����F�� UךU���u�u�u�u�w�}��������A��V�����:�!�:�
��8�(��O���T��Q1�����3�
�d�
�'�/����&��ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z���
������T��[���_�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���m�3�8�b�w�3�W���Qۇ��P	��C1�����e�h�2�%�1�m���&����^��G1�����|�u�=�;�w�}�W���Y���F��d1�����0�8�&�;�8��;���H˹��T9��X��Hʲ�%�3�e�3�f����A����A��E ��N���u�u�u�u�w�}�Wϸ�&����l��Z1�������<�d��8�(��K���T��Q1����
� �c�m�6���������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�m�3�8�f�t�^Ϫ����F�N��U���u�3�
�����������P��S����� �c�d�%�l�}�W���Y���F������,� �
�
�2��@��E�ƫ�C9��hX�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�F������F��SN��´�
�<�
�1��k�^�������F�N��U���u�u�3�
���E�������9��P1�F���h�3�
���o�8���Kù��U��]��F�ߊu�u�u�u�w�}�W���*����2��x��Gڊ�
�0�
�c�c�a�W���������C1�*ي� �d�`�
�d�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�|�!�0�]�}�W���Y���F�Q=��8���g��!�b�f�/���N��� ��O#��!ػ� �
�
�
�"�l�E݁�J���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���d�3�8�d�~�t����s���F�N��U���3�
���.�(�(�������lW��1����m�u�h�2�'�;�(��&����F�N��U���u�u�3�
������&����Z��hX��*���
�c�m�i�w�/�(���N�ѓ�]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��F���PӒ��]l�N��U���u�u�u�'�0�j�@��Y����U��Y��G�ߊu�u�u�u�w�}�W�������F�	��*���c�d�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y���R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����G^��D��\ʴ�1�;�!�}�'�>��������lV�	��*���
�
�e�3��j�(�������O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��ӊ�&�
�|�u�%�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O��Y
�����4�
�:�&��2����Y�ƫ�C9��1��F���
�d�
�%�3�3�^������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�u�=�;�w�}�W���Y���F��R	��A���h�2�%�3��m�(��s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�b�u�9�}��������]��[����h�2�%�3�g�;�F߁�����l��S��\���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�l�1�0�O������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���4�1�;�!��-��������Z��S�����
�
�
�
�"�k�O���&����O�N���ߊu�u�u�u�w�}�W�������F�	��*���b�g�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y���R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����G_��D��\���'�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�`�1�0�F�������\�V�����
�:�<�
�w�}����&ù�� 9��hX�*���1�;�|�|�~�)��ԜY���F�N��Uʧ�2�b�b�i�w�/�(���N�ѓ�]ǻN��U���u�u�u�u�2��A���DӁ��l �� \����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C�����;�%�:�0�$�}�Z���YӖ��P��F��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y�����Yd��U���u�u�u�<�w�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����
O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�e�~�t����s���F�N��U���'�2�b�b�k�}��������l��=N��U���u�u�u�u�w�8�(��Y����A��B1�G���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���u�0�!�&�6�8�_���7����^O��QN��ʦ�4�0�8�6�>�8�W��Y����C9��h��*���<�;�%�:�w�}����
����C9��h��Yʴ�
�0�u�'���(���I����Q��V�����u�'�
�
���(���O�ޓ�C9��Y����<�
�1�
�a�q�����֓�lW��Q��Cۊ�%�1�;�|�w�}�������F���ʴ�
��3�8�>�W�W���Y���F��R �����
�!�
�&��}�I�ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�%�$�:����O���F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�;���s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���g�3�8�d�j�}�W���Y���F�N�����
�&�u�h�6��#���J����lT��N��U���u�u�"�0�w�-�$�������^9��
P��U���u�u�u�u�w�}����*����Z�V��!���a�3�8�f�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N������3�8�i�w�-�$���ƹ��^9��=N��U���u�u�u�=�9�<�(���
�ӓ�@��S����u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y�����YN��*���&�c�3�8�b�`�W���Y���F�N��U����
�&�u�j�<�(���
�ѓ�@��d��U���u�u�u�"�2�}����&����U��N��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�m�3�8�`�W�W���Y���F��R �����
�!�
�&��}�I�ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�4��2��������F�P�����3�d�
� �a�e�������O��_��U���u�u�u�u�w�}�W�������l ��R������&�l�3�:�e�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N������3�8�i�w�-�$����֓�@��d��U���u�u�u�"�2�}����&����l ��hW��K�ߊu�u�u�u�w�}�W���	����U��S�����
�!�d�3�:�l�L���Y���F���ʴ�
��&�d��.�(��D��ƹF�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�d�h�u�w�}�W���Y���F��G1��*���u�h�4�
��.�F܁�
����l�N��U���u�"�0�u�'��(���J����lW��
P��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�d�W�W���Y���F��R �����
�!�a�3�:�l�W���s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}�6�����&����P9��
N�����e�3�d�
�"�k�F���&����O������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d��.�(��s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���������� ]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!�b�;���Y���F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u��������_	��T1�Hʲ�%�3�e�3�d�;�(��&����\��G�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�k����H��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���Hƹ��^9��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���;�4�
��$�l�(���&���FǻN��U���u�u�u�u�'��(���Y����C9��h��B���8�d�n�u�w�}�W���Yӑ��]F��h=����
�&�
�c�j�}�W���Y���F�N�����
�&�u�h�6��#���H˹��^9��d��U���u�u�u�"�2�}����&����l ��h_�H���u�u�u�u�w�}�W�������l ��R������&�d�
�$��O�ԜY���F�N�����%��
�!�n�;���Y���F�N��U���u�u�4�
��;���Y����g9��^�����l�_�u�u�w�}�W�������C9��h��E���8�d�u�k�]�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�=�;�6��#���K¹��^9��S����u�u�u�u�w�}�W���7����^F���&���!�g�3�8�e�f�W���Y���F��_������&�g�
�$��F��Y���F�N��U���u�%��
�$�}�JϿ�&����GW��D��N���u�u�u�u�w�*��������[�d��U���u�u�u�u�w�<�(������F��o6��-���������/��Y���F��Y
�����_�u�u�;�w�/����B���F������u�&�<�;�'�2����Y��ƹF��G1�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�E݁�
����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���K����lT��G�����_�u�u�u�w�}�W�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�:�2�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������]F��X�����x�u�u�4��9����
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�|�u�w�?����Y���F��QN�����}�%�6�;�#�1����H����C9��V��\ʴ�1�}�%�6�9�)���������D�����
��&�d�1�0�G���Y����l�N��U���u�4�
�1�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���'�4�,�4�$�:�W�������K��N�����0�1�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��_��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���u�=�;�_�w�}�W���Y�ƭ�l��S��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-���� ���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��S1�G���&�<�;�%�8�8����T�����D�����d�g�
�&�>�3����Y�Ƽ�\��DF��*���3�8�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��m�@��Yۇ��P	��C1��D��h�4�
��1�0�E�������T��UךU���;�u�'�6�$�f�}���Y���R��^	�����e�b�4�&�0�}����
���l�N��*���
�1�
�e�`�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���J���N��h�����#�
�u�u�'��(���Q�ƨ�D��_��N���u�0�1�%�8�8��Զs���K��G1�����1�d�a�u�$�4�Ϯ�����F�=N��U���&�2�7�1�f�i�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&����Z������!�9�d�d�j�<�(��������Y��A���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�e�f�<����Y����V��C�U���4�
�<�
�3��G�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������S��S�����:�&�
�#��}�W���:����^N��
�����d�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�l�@Ͽ�
����C��R��U���u�u�4�
�>�����IĹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ہ�����p	��E�����4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�F��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�4� �;�2����&����R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�d�c�4�$�:�W�������K��N�����<�
�1�
�f���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�6�(��������V9��V�����u�u�7�2�9�}�W���Y���F������7�1�d�c�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hZ�����9�:�!�:���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�@ʴ�&�2�u�'�4�.�Y��s���R��^	�����g�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ފ�4� �9�:�#�2�(���&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��D���i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ғ�R��[-�����
�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Z�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lR��V �����!�:�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����U��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�i�:�������G��h��*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��C���
������T��[���_�u�u�%�$�:����H�Փ�@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q����4����_%��C��*���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�a��;�6���������l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�`�u�$�4�Ϯ�����F�=N��U���&�2�7�1�f�o��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�a��3��������l��h�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�`�w�`�_���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��8���4��;�'�;�8�A���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��@��4�&�2�u�%�>���T���F��h��*���
�`�m�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�E���D�έ�l��D��ۊ�u�u�%���.�_�������S�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����d�4�&�2�w�/����W���F�V�����1�
�c�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�4� �;�2����&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����d�d�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lR��V �����!�:�
�
��-����P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Bڊ�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��h[�����
�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�`��3����I����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����b�u�&�<�9�-����
���9F������7�1�d�l�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�`��;�2�8�F���&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����V9��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�f�e�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(�������9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�m�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h<�����
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��l4��P��*ي�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��N���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�`��;�0�2�n�������9F���U���6�&�n�_�w�}�Z���	����l��h\�U���<�;�%�:�2�.�W��Y����C9��P1����c�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��@���;�0�0�a�6�����Y����V��=N��U���u�u�u�u�w�-��������P�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u������&����R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�g�`�4�$�:�W�������K��N�����<�
�1�
�f���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�6�:�(���&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��G���i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ӓ�R��h��*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��E���
������T��[���_�u�u�%�$�:����K�ғ�@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q����+����l��h�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�g�w�`�_���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��'���0�0�c�4��1�^��Y����]��E����_�u�u�x�w�-�������� U��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��]�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��e�����b�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���J�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�4�0��(؁�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��G��4�&�2�u�%�>���T���F��h��*���
�a�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1�U���
�4�2�
���������F��P��U���u�u�u�u�w�}��������W9��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�B�������l^��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�`�w�.����	����@�CךU���%�&�2�7�3�o�F���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�b������ߓ�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����`�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��Y	�����4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���IӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&Ź��A��C��*���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�c��'�:�)����&ù��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����g�l�4�&�0�}����
���l�N��*���
�1�
�c��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�4�6�8�����ד�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����c�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��E�����
�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Y�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lQ��V��*���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�b��<�$�8�G���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��E���&�<�;�%�8�8����T�����D�����f�c�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^�����<�&�0�f�<�(���P�����^ ךU���u�u�u�u�w�}��������lU��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������9��h��\��u�u�0�1�'�2����s���F������7�1�f�`�6�.��������@H�d��Uʴ�
�<�
�1��l�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��<����&����l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����`�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l!��Y��*؊�%�#�1�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ϯ�N����]��h]�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�e�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��B���<�&�0�f�6�����B����������n�_�u�u�z�}��������lU�������%�:�0�&�w�p�W�������T9��S1�F���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F�� 1�����0�a�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����J���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�6�3�(���&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����g�4�&�2�w�/����W���F�V�����1�
�a�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�4�;���(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Z�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����>����l��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�b�}����Ӗ��P��N����u�%�&�2�5�9�D�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�j�0���
����l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�`�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��p�����c�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����J����@��YN�����&�u�x�u�w�<�(���&���� P��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����t��D1��B���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�n�G��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�4�;�
����������F�R �����0�&�_�_�w�}�ZϿ�&����Q��X����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���;�
�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������
F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�`������ޓ�C9��SG����u�;�u�'�4�.�L�ԶY���F��h��*���
�b�u�&�>�3�������KǻN�����2�7�1�f�o�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��B���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��Z��R1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�n�W�������A	��D�X�ߊu�u�%�&�0�?���&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&���� ^�
N�����
�&�}�u�8�3���Y�ƭ�l��D��ۊ�|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�o�}����Ӗ��P��N����u�%�&�2�5�9�D�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�d�$�������lV��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����&�0�e�4��1�^��Y����]��E����_�u�u�x�w�-��������
P��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��W�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��d�����0�d�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����J���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�>�3����&¹��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����a�`�4�&�0�}����
���l�N��*���
�1�
�e��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�e��#�2�����֓�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����e�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�V��R�����
�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6��������� F��D��U���6�&�{�x�]�}�W���
����W��]�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lW��~ �����
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����K���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�d�
�9�(����I����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����f�u�&�<�9�-����
���9F������7�1�a�g�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�d�
�;�"�.��������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��F���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&�ד�]��D1��D���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���H����F��R1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�c�l�K��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*����%�!�
����������F�R �����0�&�_�_�w�}�ZϿ�&����Q��[����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*���
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����D���%�!�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����S��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�l�(�������lU��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�`�w�.����	����@�CךU���%�&�2�7�3�i�N���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�f�����
����l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�`�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��h'�� ���0�a�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�W��Y�����`�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���A�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�d��'�)�(���&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����b�4�&�2�w�/����W���F�V�����1�
�b�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�d��%�#��(ف�	����l�N�����u�u�u�u�w�}�W�������T9��S1�B��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�H¹��C��h��*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��O���
������T��[���_�u�u�%�$�:����M�ޓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��V��H���%�6�;�!�;�l�F������l ��]�����:�f�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��N���
������T��[���_�u�u�%�$�:����M�ѓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��Y��H���%�6�;�!�;�l�F������l ��X�����:�c�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��G���
������T��[���_�u�u�%�$�:����L�Г�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��X��H���%�6�;�!�;�l�F������l ��_����!�u�d�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h[�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�b�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h[�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�m�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h[�U��}�%�6�;�#�1�F��DӇ��p5��D��Aʱ�"�!�u�a�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����L�ƭ�@�������{�x�_�u�w�-��������U��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��@���h�}�%�6�9�)����H����C9��h��]��1�"�!�u�o�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lS��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����u�:�;�:�n�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lS��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����e�1�"�!�w�m�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��X�����;�%�:�u�w�/����Q����G��N��A���;�4��;�%�1��������W9��h��Yʥ�a��;�4��3�����ד�C9��S1��*���y�%�a��9�<�4�������lT��G1�����
�<�y�%�c�����:����\
��h]�����1�<�
�<�{�-�C�������\��X��*ފ�%�#�1�<��4�[Ϯ�M����F��X �����
�
�%�#�3�4�(���UӖ��l+��B�����:�
�
�
�'�+����&������h#�� ���:�!�:�
����������@����*���2�
�
�
�'�+����&������h<�����
�
�%�#�3�4�(���UӖ��l4��P��*؊�%�#�1�<��4�[Ϯ�L����T��h]�����1�<�
�<�{�-�B�������lR��G1�����
�<�y�%�b������ӓ�C9��S1��*���y�%�`��9�8��������W9��h��Yʥ�`��;�0�2�j��������l��N��@���;�0�0�m�6���������F��1�����0�l�4�
�;������Ƽ�9��E�����
�
�
�%�!�9��������lP��V�����&�0�d�4��1�(���
���C9��p�����e�4�
�9��3����Y����t��D1��D���
�9�
�;�$�:�W���&����@9��1��*���
�;�&�2�w��(������� 9��h��*���&�2�u�
��<����&ǹ��l��h�����u�
�
�4�9��(ځ�	����l��D��U���
�4�;�
����������@����*���;�
�
�
�'�+����&������h)�����
�
�%�#�3�4�(���UӖ��l!��Y��*ӊ�%�#�1�<��4�[Ϯ�@����]��h��*���#�1�<�
�>�q����*����_��h_�����1�<�
�<�{�-�F߁�����]��R1�����9�
�;�&�0�}�(���0����@9��1��*���
�;�&�2�w��F���	����V9��V�����;�&�2�u��l�>�������9��h��*���&�2�u�
�f�����&����R��[
�����2�u�
�d��-����&ǹ��l��h�����u�
�d��'�)�(���&����_��Y1�����
�d��%�#��(ف�	����l��D�����u�0�<�_�w�}�W���Y���F��h��*���
�c�u�h��-�Fށ�����l��h�����<�
�<�u�w�-��������Z��N��U¥�d�
�;� �$�8�B���&����Z��^	��U���6�;�!�9�0�>�G����μ�W��Y�����a�4�
�9��3����DӇ��P	��C1�����e�u�'�}��l�>������� 9��h��*���&�2�h�4��2��������O��EN��*����%�!�
����������@��
N��*���&�
�:�<��t����	����z��C��*ۊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�d��3�����֓�C9��S1��*���u�u�%�6�9�)�������\�G1�*���%�<�!�
����������@��
N��*���&�
�:�<��t����	�ߓ�Z��[��*ۊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�l��:�����֓�C9��S1��*���u�u�%�6�9�)�������\�G1��2���&�0�l�4��1�(���
�����T�����2�6�e�u�%�u�(؁�����V9��V�����;�&�2�h�6�����&����P9����]���
�4�;�
����������@��
N��*���&�
�:�<��t����	�ѓ�R��h��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�b��>�.��������W9��h��U���%�6�;�!�;�:���Y���C9��p�����a�4�
�9��3����DӇ��P	��C1�����e�u�'�}������&����R��[
�����2�h�4�
�8�.�(�������	����*���;�
�
�
�'�+����&����F��h�����:�<�
�|�8�}����>����l��h�����<�
�<�u�w�-��������Z��N��U¥�b��<�&�2�m��������l��S�����;�!�9�2�4�m�W���Q����c��Z�����
�
�%�#�3�4�(���Y�ƭ�l��D�����
�|�:�u�'�k�'�������@9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�4�2���(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l4��P��*Ҋ�%�#�1�<��4�W���	����@��X	��*���:�u�%�`��3����N����E
��^ �����u�%�6�;�#�1����I�ƣ�N��1�����0�c�4�
�;���������C9��Y�����6�e�u�'���(�������9��h��*���&�2�h�4��2��������O��EN��*ߊ�4�2�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�L����T��h]�����1�<�
�<�w�}��������\��h^�����%�`��;�2�8�E���&����Z��^	��U���6�;�!�9�0�>�G����μ�9��Y	�����4�
�9�
�9�.�������]��[����u�'�}�
��<����&ù��l��h�����h�4�
�:�$�����&����AF��hZ�����9�:�!�:���(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l+��B�����:�
�
�
�'�+����&����F��h�����:�<�
�|�8�}����4����_%��C��*���
�%�#�1�>�����Y����\��h�����|�:�u�%�c�����:����\
��hZ�����1�<�
�<�w�}��������\��h^�����%�a��;�6���������l��A�����<�u�u�%�4�3��������F��F��A���;�4��;�%�1��������W9��h��U���%�6�;�!�;�:���Y���C9��z�����;�'�9�0�f�<�(���&����Z������!�9�2�6�g�}����&ǹ��]��t�����0�e�4�
�;���������C9��Y�����6�e�u�'��-��������C9��Y�����6�e�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��A���
������T��[���_�u�u�%�$�:����N�Г�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��X��H���%�6�;�!�;�l�F������l ��_����!�u�f�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��hV�U��}�%�6�;�#�1�F��DӇ��p5��D��Bʱ�"�!�u�b�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����H�ƭ�@�������{�x�_�u�w�-��������S��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��D���h�}�%�6�9�)����H����C9��h��]��1�"�!�u�n�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������l^��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����g�1�"�!�w�o�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����������^	�����0�&�u�x�w�}��������W9��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��l+��B�����:�
�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������Z�F��*���&�
�:�<��}�W���&����R
��Y�����e�4�
�9�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�n�u�u�2�9��������9l�N�U���&�2�6�0��	���&����
F��D��U���6�&�{�x�]�}�W���
����@��d:�����3�8�l�4�$�:�(�������A	��D�����2�7�1�`�g�W�W�������F�N�����4�
�<�
�3��@�������9F�N��U���u�%�&�2�4�8�(���
����U��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��^�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���H¹��^9�������%�:�0�&�w�p�W�������T9��R��!���d�
�&�
�g�<����&����\��E�����%�&�2�7�3�h�O�ԜY�Ʈ�T��N��U���<�u�4�
�>�����N����[��=N��U���u�u�u�%�$�:����&����GW��Q��D���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GW��Q��D���&�<�;�%�8�8����T�����D�����
��&�d��.�(�������]9��X��U���6�&�}�%�$�:����L���F�U�����u�u�u�<�w�<�(���&����V�����ߊu�u�u�u�w�}��������B9��h��G���8�d�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�g�3�:�l�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��F���8�d�u�&�>�3�������KǻN�����2�6�0�
��.�F܁�
����l��^	�����u�u�'�6�$�u��������l^��d��Uʷ�2�;�u�u�w�}��������T9��S1�D���=�;�_�u�w�}�W���Y����Z��D��&���!�f�3�8�f�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�n����H�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�a�3�8�f�}����Ӗ��P��N����u�%�&�2�4�8�(���
����U��]�����;�%�:�u�w�/����Q����Z��S
��C���u�u�7�2�9�}�W���Yӏ����D�����b�c�u�=�9�W�W���Y���F��h��*���$��
�!�c�;���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���M����lW��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!�b�;���Y����T��E�����x�_�u�u�'�.��������l��1����
�&�<�;�'�2�W�������@N��h��*���
�a�|�u�w�?����Y���F��QN�����2�7�1�`�g�}����s���F�N�����<�
�&�$����������F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����S��D��A��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$����������F��D��U���6�&�{�x�]�}�W���
����@��d:�����3�8�d�
�$�4��������C��R�����<�
�1�
�g�l�}���Y����]l�N��Uʼ�u�4�
�<��9�(��H�Ƹ�V�N��U���u�u�4�
�>�����*����P��D��@��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��D܊�&�
�`�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�>�����*����^��D��Bʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�m�1�0�F؁�
����l��TN����0�&�4�
�>�����I��ƹF��R	�����u�u�u�3��-��������T�C��U���u�u�u�u�w�<�(���&����l5��D�*���
�b�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��j�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�*���
�m�4�&�0�}����
���l�N��*���
�&�$���)�N�������R��P �����o�%�:�0�$�<�(���&����S��=N��U���<�_�u�u�w�}����	����l��h[�\ʡ�0�u�u�u�w�}�W�������T9��R��!���d�
�&�
�o�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�f�����A���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���d�3�8�e�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&����9��D��*���6�o�%�:�2�.��������W9��d��Uʷ�2�;�u�u�w�}��������T9��S1�\ʡ�0�u�u�u�w�}�W�������T9��R��!���d�3�8�e�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�d�1�0�G��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��Gڊ�&�
�l�4�$�:�W�������K��N�����<�
�&�$����������
9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��D���!�0�u�u�w�}�W���YӇ��@��T��*���&�g�
�&��d�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�o�(���&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�g�
�&��l�����Ƽ�\��D@��X���u�4�
�<��.����&����l ��h\�����2�
�'�6�m�-����
ۇ��@��U
��D��|�u�u�7�0�3�W���Y����UF��G1�����1�d�g�|�#�8�W���Y���F������6�0�
��$�o�(���&���F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
����U��_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�o����HӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����d�f�|�u�w�?����Y���F��QN�����2�7�1�d�d�t����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l ��h_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�i����JӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����a�m�_�u�w�8��ԜY���F��F��*���
�1�
�m�~�)����Y���F�N�����2�6�0�
��.�C������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
�ғ�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�b�;�������]F��X�����x�u�u�4��4�(�������@��Q��A���&�2�
�'�4�g��������C9��P1����a�|�u�u�5�:����Y����������7�1�d�a�~�)����Y���F�N�����2�6�0�
��.�B������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
�ӓ�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�a�;�������]F��X�����x�u�u�4��4�(�������@��Q��@���&�2�
�'�4�g��������C9��P1����g�|�u�u�5�:����Y����������7�1�d�g�~�)����Y���F�N�����2�6�0�
��.�A������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
�Г�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�`�;�������]F��X�����x�u�u�4��4�(�������@��Q��C���&�2�
�'�4�g��������C9��P1����b�_�u�u�2�4�}���Y���Z �V�����1�
�l�|�#�8�W���Y���F������6�0�
��$�j����O���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���N����lP�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�m�1�0�@Ͽ�
����C��R��U���u�u�4�
�>�����*����9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��@��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�d�|�!�2�}�W���Y���F��G1�����0�
��&�o�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�l�3�:�e�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�D�ߊu�u�0�<�]�}�W���Y���R��^	�����f�|�!�0�w�}�W���Y�����D�����
��&�l�1�0�O��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�N������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�Wϸ�&����|��^�� ��f�
�d�i�w��9���6����9��P1�����a�f�%�n�w�}����<����G9��h ��*��� �d�f�
�e�a�WǸ�&����|��^�����!�<�3�
�c�d�����ƭ�l��D�����m�e�e�e�~�W�W���*����K)��h_�����;�
�
� �f�o�(��E�ƾ�T9��UךU����-� ��9�(�(���H����
P��G]��H�ߊu�u�u�u��%�"�������V��B1�D���u�=�;�}�2���������
S��G\��\��r�r�u�9�2�W�W���Y�Ƽ�W��Y�����e�<�
�<�l�}�Wϸ�&����gT��B��E���3�
�d�d�'�}�JϮ�+����G9��h��D��
�`�_�u�w�����-����G9��h]�� ��`�
�f�i�w�}�W���YӀ��K+��c\�� ���e�g�3�
�f�l�������@��C��*���3�
�d�b�'�u�^��^���V
��d��U���u�%�d�
�9�(����J����@��=N��U���-� ��;�"��G���&����CW�
N��'���9�
�m�3��o�(��s���U5��z;��G���!�g�
�;�2�-�!�������
9��R�����9�2�6�#�4�2�_���������R����
� �m�d�'�t�\ϫ�
����WN��h�����#�m�d�|�]�}�W���������C1�*���0�%��f�1��G���	�����h�����0�!�'� �$�:����&����_��1��*��d�%�|�~�"�.����Q����\��h��M��|�_�u�u��%�"�������V��Y1��!���
�
� �d�c��D��Y���F���*؊�
�
�l�6�$���������S��N�����&�9�!�%��i����I�ѓ�N��S��D���0�&�u�u�w�}�Wϭ�����l��Q��E���%�n�u�u�1��:���K����lT��^ �����0�3�
�`��n�K���Y���F��R��*���
�
�4�!�4�.�(���A�ӓ� F��R �����!�%�
�
�"�e�@���Q���A��N�����u�u�u�u�$�1��������U��G]�U���3�
���e�����H����R��h�I���u�u�u�u�1��:���K����lQ��B1�Eڊ�d�"�0�u�$�1����&�ԓ�F9��X��G��u�u�d�|�2�.�W���Y��� ��O=�����
�
�0�
�`�k�}���Y����~3�� �����3�
�a�e�'�}�JϮ�+����G9��h��D��
�`�_�u�w�����-����G9��^ �����
�
� �d�e��E��Y����_	��T1�����}�;�<�;�3�-�%�������U��\�����~� �&�2�2�u��������EW��(��3���_�u�u��/��#ݰ�����Z��G:�����
�f�g�%�w�`�}���Y���A��1�����d�6�&�
�6�)����K�ғ� F��R �����!�%�
�`�1��D���	����[�I�����u�u�u�u�w�.����	����U��W����_�u�u�x�0�-��������U�� V�����u�&�<�;�'�2����Y��ƹF��E��*ڊ�
�e�3�
�`�����&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:��݊�&�
�y�4��4�(�������@��Q��B�ߊu�u�0�<�]�}�W���Y���N��h�����:�<�
�u�w�-���������T�����2�6�d�h�6�����
����g9�� 1����u�'�}�%�4�3��������[��G1�����0�
��&�o�;���P����[��=N��U���u�u�u�'���(���I����Q��V����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}�����֓�lW��Q��BҊ�%�6�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���'�
�
�
��m����N˹��l��E��Hʲ�%�3�e�3�f����A����@��C1��*���'�
�0�n�w�}�����֓�lW��Q��BҊ�;�-�e�i�w�1�1���;����F��C1�*���
�0�
�c�n�W�W���T�ƫ�C9��1��Dۊ� �c�d�4��8�����Ƽ�\��D@��X���u�2�%�3�g�;�Fށ�����l��T�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�f�����J�ƭ�l��h�����
�!�f�3�:�l�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�4�
�8�.�(�������F��h��*���$��
�!�c�;���PӉ����T�����2�6�d�h�6�����
����g9��]�����g�|�|�!�2�}�W���Y���F��E��*ڊ�
�d�3�
�a�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʲ�%�3�e�3�f����H����P�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӁ��l ��h��D���
�c�
�%�$�<���Y����U9��Q1�*���c�d�4�
�#�/�(���
����l��d��Uʲ�%�3�e�3�f����H����t��r������0�
�`�k�}�(ف�����G��h��*���&�2�_�u�w�/�(���&����l ��X������2�<�&�o�8�G��Y����t��D1��E���
�<�n�u�w�:����I����9��hX�*�����4�;���(���DӖ��l!��Y��*ۊ�;�&�2�_�w�}����&ù��W��B1�D���
��'�;�2�d���E�Ƽ�9��Y	�����<�
�<�n�w�}�����֓�lW��Q��Cۊ�;���4�0��(���Y����lS��V ��*���
�;�&�2�]�}�W���&����U9��h��C���<�
�!�!���(���Y����_9��r*��6���!� �
�b�2�m����H����9F�	��*���
�
�d�3��k�(���/����[��R	��F��u�u�2�%�1�m���&����W��Y1��*���h�%�c��%�0����&����Z��^	�U���2�%�3�e�1�l�(���O�ד�]9��D��A��u�
�
�<�9�1�(���&����Z��=N��U���2�%�3�e�1�n����H˹��l��V�����'�6�&�{�z�W�W�������9��1��*��
�%�6�
�$�4��������C��R�����0�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���M����lW��	��*���
�
�d�3��k�(�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������_	��T1�Hʴ�
�<�
�&�&��(���L����lW����]´�
�:�&�
�8�4�(���Y����Z��D��&���!�a�3�8�f�t�������R��X ��*���<�
�u�u�%��(߁�&�ד�F9��1��*���0�|�|�|�#�8�W���Y���F�	��*���
�
�
� �a�e�������R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���'�
�
�
�����A����P�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӁ��l ��h��*���c�m�4�
�#�/�W������lV��h]�� ��m�4�
�!�%���������V��N�����3�e�3�f�1��Fׁ�����]��h��U��%�b��<�$�8�E���&����9F�	��*���
�
�
� �a�e��������9��N�U���
�4�;�
���������F��G1��E���f�3�
�d��3�0���
�ғ�lT�
N��B���<�&�0�a�>����Y����A��h^��*ي� �c�m�<��<����&����[��hY�����
�
�
�;�$�:�}���Y����U9��Q1�����d�
�;��>�.�C���M���C9��p�����c�<�
�<�l�}�WϹ�	����l ��h��C���<�
�4�;���(���DӖ��l!��Y��*݊�;�&�2�_�w�}����&ù�� 9��hX�*����<�&�a�2�k�K���&Ĺ��Z��R1�����<�n�u�u�0�-�����Փ�F9��1��*���;�
�
�
�w�`����>����l��h�����_�u�u�'���(���&����^��Y1������;�'�9�f��(���DӖ��l+��B�����:�
�
�
�9�.��ԜY�ƫ�C9��1��F���
�d�
�;��3��������lW��R1�I���
�
�4� �;�2����&����Z��^	�U���2�%�3�e�1�n����H˹��l+��B�����:�
�g�0�e�a�W���&����R
��Y�����g�<�
�<�l�}�WϹ�	����l ��h��C���<�
�4� �;�2����&�ԓ�lU�
N��A���;�4��;�%�1��������T]ǻN�����
�
�
�
�"�k�O���&����R
��Y����
�
�u�h�'�i�:�������G��h��*���&�2�_�u�w�/�(���&����U��V�����;�4��;�%�1�F݁�&�����h#�� ���:�!�:�
���������F��G1��E���f�3�
�d��3�:�������G��h_����i�u�
�
�6�(��������V9��^ ����u�u�2�%�1�m��������9��h#�� ���:�!�:�
�e�8�@��Y����~��V�����9�0�b�<��4�L���YӁ��l ��h��*���c�m�<�
��o���E�ƪ�l��R1�����=�0��4�2��(���&����Q��d��Uʲ�%�3�e�3�d�;�(��&����e9��R1�I���
�d��%�#��(ف�����l�N�����e�3�f�3��l�(���)����V9��S��&����,� �
�f�l����H����9F�	��*���
�
�
� �a�e����/�ԓ�lU�
N��*�����!��5�/����A�ד�V��W����u�'�
�
���(���O�ޓ�]9��Y	��B���e�i�u�
��<����&����l��d��Uʲ�%�3�e�3�d�;�(��&����R��hY��*���h�%�`��9�8��������T]ǻN�����
�
�
�
�"�k�O���&����V9��R1�I���
�
�4�2���(���
����F�P�����3�f�3�
�f���������l��R������;�0�0�b�4�(���B�����h��*���
� �c�m�>�����&Ĺ��F���*���2�
�
�
�9�.��ԜY�ƫ�C9��1��F���
�d�
�;��3�������F��1�����0�b�<�
�>�f�W�������lV��h]�� ��m�<�
�4�0��(���Y����lS��V ��*���
�;�&�2�]�}�W���&����U9��Q��DҊ�;��;�0�`�8�@��Y����a��R1��L���
�<�n�u�w�:����I����l ��_������d�0�e�k�}�(ف�����G��h��*���&�2�_�u�w�/�(���&����U��V�����
�
�
�u�j�-�F߁�����]��R1�����<�n�u�u�0�-�����Փ�F9��1��*���0�
�u�h�'�d�$�������lW��Y1���ߠu�u�x�u�%����N����R��P �����&�{�x�_�w�}��������l��V�����'�6�o�%�8�8�ǿ�&����P��h=�����3�8�e�u�'�>�[Ͽ�&����P��h=�����3�8�b�u�'�.��������l��h��*���4�
�<�
�$�,�$����ӓ�@��B�����2�6�0�
��.�Fց�
����F��h��*���$��
�!�c�;���UӁ��l ��h��D���
�c�
�%�3�3�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y����\�V�����
�:�<�
�w�}����P�ƣ�N��h�����:�<�
�u�w�-��������`2��CV�����|�:�u�4��2��������F�V�����&�$��
�#�����PӉ����T�����2�6�d�h�6�����
����g9��[�����a�u�'�}�'�>��������lW������6�0�
��$�l�(���&���\������!�9�2�6�f�`��������V��c1��Dފ�&�
�f�u�9�}��������_	��T1�Hʲ�%�3�e�3�f����H����W	��G��U���;�_�u�u�w�}�W�������lP��h��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�:����&����P�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h��C���:�6�1�u�$�4�Ϯ�����F�=N��U���
� �c�b�8�>����
����l��TN����0�&�4�
�>�����*����T��D��D���%�&�2�6�2��#���Hù��^9�������6�0�
��$�o�(���&���R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�a�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF������!�9�2�6�f�`��������V��c1��Gڊ�&�
�l�u�%�u��������\��h_��U���&�2�6�0��	��������F��F��*���&�
�:�<��}�W���
����@��d:��ߊ�&�
�|�:�w�<�(���
����T��N�����<�
�&�$����������O����ߊu�u�u�u�w�}��������l	��X
��I���%�6�;�!�;�o�F�ԜY���F��D��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��l�W���Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����U��Y�����0�i�u�%�4�3����K����F�N�����u�u�u�u�w�}�WϹ�	����^��X�����h�w��n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӁ��l ��V�����&�<�;�%�8�8����T�����h��C���%�
�&�<�9�-����Y����V��G1�*��� �&�0�d�>��������T9��R��!���d�
�&�
�f�}����M����V��Y����<�
�&�$����������F��h��9����!�g�
��8�(��@�ƪ�l��{:�� ��� �!�%�,�a�l����H������D�����
��&�g��.�(��Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����a�u�%�&�0�>����-����9��Z1�\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���T��Q��M݊�e�i�u�0��i�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�f�t����Y���F�N��U���
� �c�b�'�}�Jϸ�&����g��C1�����9�
�
�
�2��A��s���F�R�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����P��D��@���u�=�;�_�w�}�W���Y�ƫ�C9��hX�*��i�u�0�
�b�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�a�|�#�8�W���Y���F�	��*���c�b�%�u�j�-�Fށ�����l��h�����_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����l ��h_��U���;�_�u�u�w�}�W�������lP��h�I����-� ��9�(�(���H����lW��UךU���u�u�9�0�]�}�W���Y���T��Q��M݊�e�i�u����/���!����k>��o6��-������n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӁ��l ��V�����&�<�;�%�8�8����T�����h��C���%�
�&�<�9�-����Y����V��G1�*��� �&�0�d�>����	����z��C��*؊�;�&�2�u�'�.��������l��1����y�'�2�b�e�}����O����C9��P1������&�d�
�$��[ϸ�&����gT��B��*ۊ�0�
�b�e�w�-��������`2��C\�����d�y�4�
�>�����*����9��Z1�U���&�2�6�0��	��������F��h��*���$��
�!�a�;���P�����^ ךU���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�G�������F��R ��U���u�u�u�u�0�-����AĹ��Z�Q=��8���g��!�b�f�/���N��ƹF�N�����u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u�'�
�"�k�@���Y����V��Y�U���u�u�0�&�1�u�_�������l
��^��U���%�&�2�6�2��#���Hù��^9����]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�b�t�W������F�N��Uʲ�%�3�
�m��l�K�������]ǻN��U���9�<�u�}�'�>��������lW������6�0�
��$�h����M����[��=N��U���u�u�u�'��(�A���	�����1�����
�
�
�;�$�:�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����
�m�
�d�k�}�(���0����@9��1��*���n�u�u�u�w�8����Y���F�N����� �c�b�%�w�`�U���!����k>��o6��-���������U�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�P�����l�
�0�4�$�:�W�������K��N�����3�
�l�
�2�<����&����\��E�����%�&�2�6�2��#���H����lV�V�����%�&�2�6�2��#���A����lQ�V�����&�$��
�#�����UӇ��@��T��*���&�d�
�&��i�W���
����@��d:�����3�8�d�y�6�����
����g9��Z�����f�u�'�
���(�������9��h
���ߊu�u�0�<�]�}�W���Y���N��h�����:�<�
�u�w�-��������`2��C_�����|�:�u�:��<�(���
����T��N�����0�|�:�u�6�����&����P9��
N��*���
�&�$���)�(���&����AF��G1�����9�2�6�d�j�<�(���&����l5��D�����m�u�'�}�'�>��������lW������6�0�
��$�l�(���&���\�V�����
�:�<�
�w�}��������B9��h��L���8�d�|�:�w�u��������\��h_��U���&�2�6�0��	���&����U�V ��]���6�;�!�9�0�>�G������lV��h_�����c�
�%�1�9�t�^������F�N��U���2�%�3�
�n����Y����\��h�����n�u�u�u�w�8����Y���F�N����� �c�d�6�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�%����H����\��V�����'�6�&�{�z�W�W�������lP��h�����4�&�2�
�%�>�MϮ�������D�����
��&�d��.�(��Y����Z��D��&���!�e�3�8�n�}��������B9��h��E���8�d�y�4��4�(�������@��Q��D���%�&�2�6�2��#���L����lR�V�����&�$��
�#�k����H��ƹF��R	�����u�u�u�3��u��������\��h_��U���&�2�6�0��	���&����W�X�����:�&�
�:�>��W���	����l��F1��*���e�3�8�l�w�/�_�������l
��^��U���%�&�2�6�2��#���Kù��^9��N��U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���ƹ��^9��G�����_�u�u�u�w�}�W���&����
W��G����u�%�6�;�#�1�E��s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�c�3�:�l�^������F�N��U���2�%�3�
�n��������R��X ��*���
�n�u�u�w�}����Y���F�N��U���
� �c�d�8�>����D�Ĕ�]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�'�
� �a�l����
������T��[���_�u�u�'��(�A���	ù��@��h����%�:�0�&�%�:�@��Y����Z��D��&���!�g�3�8�f�q����N���R��^	������
�!�e�1�0�N�������J��d1�� ���;� �
�e�d�/���M����`9��p����
� �d�f��l�W���
����@��d:�����3�8�d�y�6�����
����g9��1����u�%�&�2�4�8�(���
�ӓ�@��N��*���
�&�$���)�A�������9F����ߊu�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���I����lW��N�����u�u�u�u�w�}��������9��R������-� �
�g�;�(��@����9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����H����[��=N��U���u�u�u�'��(�A���	�����hY�N���u�u�u�0�$�;�_���	����@��X	��*���u�%�&�2�4�8�(���
����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��h�^������F�N��U���2�%�3�
�n��G��Y����S��=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�B��������YNךU���u�u�u�u�%����H����[��R	��G��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�WϹ�	����_��G^��Hʳ�
���g��)�E߁�&����P��d��U���u�0�&�u�w�}�W���Y����A��B1�D���u�h�w����/���!����k>��o6��-�����w�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����U��_��Dʴ�&�2�u�'�4�.�Y��s���T��Q��Lۊ�d�4�&�2��/���	����@��h_��<���!�
�
�
�9�.����&�ד�]��D1��A���
�<�y�4��4�(�������@��h��*��u�0�
�c�{�<�(���&����l5��D�*���
�y�3�
������&����Z��h_��D���2�d�m�y�1��:���K����lQ��h��*��e�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�b�;���Y����Z��D��&���!�c�3�8�f�t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�e�1�0�F���Y����l�N��U���u�2�%�3��d�(��E�ƪ�l��{:��:���b�d�'�2�f�j�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�f�t����Y���F�N��U���
� �c�d�'�}�Jϸ�&����g��C1�����9�
�`�d�%�:�F��B���F������}�4�
�:�$�����&���R��^	������
�!�e�1�0�N����έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�!�0�u�w�}�W���Y����A��B1�D���u�h�'�2�`�o�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����
�l�
�d�k�}�(���0����@9��1��*���n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W�������F9��1��U��%�d�
�;�"�.��������T]ǻN��U���9�0�_�u�w�}�W���Y����U��_��D��u������/���!����k>��o6��-����n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϹ�	����_��T�����;�%�:�0�$�}�Z���YӁ��l ��W�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�@������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�`�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
��]���6�;�!�9�0�>�F������T9��R��!���b�3�8�c�w�/�_�������l
��^��U���%�&�2�6�2��#���L����lR�X�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�}����s���F�N�����3�
�l�
�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��E�� ��`�6�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���'�
� �c�b�-�W��	����z��C��*ފ�;�&�2�_�w�}��������l��S��*����%�!�
��������ƹF�N�����
�l�
�0�6�.��������@H�d��Uʲ�%�3�
�l��8��������\������}�%�6�y�6�����
����g9�� 1����u�%�&�2�4�8�(���
�ӓ�@��N��*���
�&�$���)�(���&��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��<�(���
����T��N�����<�
�&�$���؁�
����	�������!�9�2�6�f�`��������V��c1��@���8�a�u�'��-��������Z��S�����2�6�0�
��.�A������O��_�����u�u�u�u�w�/�(���O�ߓ�VF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��Nց����R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}��������
9��R�����b�a�_�u�w�/�(���O�ߓ�F���D���%�!�
�
��3����s���K�P�����e�
�e�4�$�:�W�������K��N�����3�
�e�
�g�<����&����\��E�����0�
�g�y�%�:�@��Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���@����lW����*��y�4�
�<��.����&����l ��hW����<�
�&�$����������J��d1�� ��� �
�d�d�%�:�F��UӀ��K'��N!��*܊�0�
�b�a�w�/�(���&����U��V�����!�'�
�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�l�3�8�f�t�W������F�N��Uʲ�%�3�
�e��m�K���*����w��C1�����d�c�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��[�����a�|�!�0�w�}�W���Y�����h��B���%�u�h�2�'�;�G���J����W��V�����;�l�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���T��Q��E݊�e�i�u�0��k�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�~�}����s���F�N�����3�
�e�
�g�a�W�������|��_��*���
�c�c�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��CW�����|�u�=�;�]�}�W���Y���T��Q��E݊�e�i�u�0��i�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���m�3�8�b�~�)����Y���F�N����� �b�b�%�w�`����N����F�N�����u�u�u�u�w�}�WϹ�	����V��G^��H���������/���!����k>��o6��-���_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������lQ��h�����2�
�'�6�m�-����
ۇ��@��T��*���&�m�3�8�`�}��������B9��h��*���
�y�4�
�>�����*����S��D��A���%�&�2�6�2��#���Hʹ��^9��N��*���
�&�$���)�G������R��^	������
�!�d�1�0�F������W��R�����:���<�f�����O���F�U�����u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����^����ߊu�u�u�u�w�}��������l��S�����;�!�9�f���3��I���F�N�����}�}�%�6�9�)���������D�����
��&�l�1�0�O����έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���:�u�4�
�8�.�(�������F��h��*���$��
�!�f�;���P����[��=N��U���u�u�u�'��(�@���	��� ��Y��*���8�&�;�:�����&����P��d��U���u�0�&�3��u��������\��h_��U���&�2�6�0��	��������F��F��*���&�
�:�<��}�W���
����@��d:�����3�8�l�|�w�5��ԜY���F�N�����
�e�
�d�k�}��������EU��(�6��n�u�u�u�w�8����Y���F�N����� �b�b�%�w�`�U���!����k>��o6��-���������U�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�P�����d�
�e�4�$�:�W�������K��N�����3�
�d�
�g�<����&����\��E�����0�
�f�y�%�:�@��Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1�Yʧ�2�b�b�u�'�.��������l��1����u�%�&�2�4�8�(���
����U��^�������!�e��(���&����F��G1��E���f�3�
�d��-��������9F����ߊu�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���L����lW��N�����u�u�u�u�w�}��������9��R�����3�e�3�f�1��Fׁ�	����F��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����V����ߊu�u�u�u�w�}��������l��S�����c�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��h��*���u�=�;�_�w�}�W���Y�ƫ�C9��hY�*��i�u��-��$����J�ד�V��X����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���@����l^����ߊu�u�u�u�w�}��������l��S�����a�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��B���!�0�u�u�w�}�W���YӁ��l �� _�����h�'�2�b�c�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��F݁�I���>��o6��-���������/���!����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�'�
� �`�o����
������T��[���_�u�u�'��(�@���	¹��@��h����%�:�0�&�6�����
����g9��1����u�%�&�2�4�8�(���
�ߓ�@��N��*���
�&�$���)�B���������D�����
��&�d��.�(������T9��R��!���d�
�&�
�g�}�$�������A��^ �����#�
�l�'�0�l�@���Y����V��=N��U���u�3�}�}�'�>��������lW������6�0�
��$�d����A�ƣ�N��h�����:�<�
�u�w�-��������`2��C_�����d�|�:�u�6�����&����P9��
N��*���
�&�$���)�F�������O��_�����u�u�u�u�w�/�(���N�ԓ�F������
�0�8�&�9�2�$�������A��X�N���u�u�u�0�$�;�_���	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��N��U´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�t�W������F�N��Uʲ�%�3�
�d��l�K���	����@��A]��F�����n�u�w�}�Wϻ�
��ƹF�N��U���'�
� �b�e�-�W��[����k>��o6��-���������/���[���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����3�
�d�
�g�<����Y����V��C�U���2�%�3�
�f��G���
����C��T�����&�}�%�&�0�>����-����l ��hV����<�
�&�$����������J��R	��@���4�
�<�
�$�,�$����ד�@��B�����b�y�2�%�1�m��������9��h�� ���m�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��Dߊ�&�
�a�|�#�8�W���Y���F�	��*���b�b�%�u�j�:����I����l ��_�����0� �;�m�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��D���8�d�|�u�?�3�}���Y���F�P�����d�
�e�i�w�8�(��B���F������}�%�6�;�#�1����H����C9��P1������&�l�3�:�e�^Ϫ���ƹF�N��U���'�
� �b�`�-�W������V��N��U���0�&�u�u�w�}�W���YӁ��l �� _�����h�w�����/���!����k>��o6��-����w�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}��������l��S��&���1�
�0�8�$�3����5����
9��P1�B��_�u�u�x�0�-����K¹����^	�����0�&�u�x�w�}��������9��h�����%�:�u�u�%�>����	����l��F1��*���
�&�
�y�6�����
����g9��[�����a�u�0�
�b�q��������V��c1��Dۊ�&�
�e�u�2��@������lV��h]�� ��m�4�
�0�"�3�O�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����M����[��=N��U���u�u�u�'��(�@���	�����h��*���
� �c�m�6���������F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!�f�;���P�Ƹ�V�N��U���u�u�2�%�1��Eށ�I���A�� Y����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���@����l^����ߊu�u�u�u�w�}��������l��S�����`�n�u�u�w�}����Y���F�N��U���
� �b�d�'�}�J���!����k>��o6��-���������/���s���F�R ����_�u�u�;�w�/����B���F��G1��*��
�d�i�u��3��������Z��D=�����m�'�2�d�a�f�W�������lW��Q��Lߊ�d�i�u�
�6�o����&����CW�N�Dʱ�"�!�u�|�]�}�W���&����l ��Y�����h�%��9��d����N¹��U��S�����f�n�u�u�;�>�!��&����S��N�U���4�g�b�
�"�d�F���Q���W��X����n�u�u�9�4��E݁�����9��R�����9�
�d�3��o�F���Q����\��XN�\�ߊu�u�:�
��n����K�ғ�F������m�
� �d�c��F��Y����W	��C��\�ߊu�u�:�
��(�@���	�����V�����
�m�
�d�d�}��������l�N��E��
�
�d�3��m�D���Y���F�N�����:�&�
�#�d�m� ���Yے��l^��Q��E���%�}�|�h�p�z�W������F�N�����g�
� �l�b�-�L���YӖ��V��1��*���d�`�
�f�k�}�W���Y����C9��Y����
�u�=�;��0�(�������P��F�U���d�|�0�&�w�}�W���Yӊ��l0��1��*��a�%�n�u�w�-�G��&¹��U��]��F��u�u�u�u�w�<�(���
����U�������8�
� �m�`�-�_���D����F��D��U���u�u�9�6��l�(���N�ӓ�]ǻN��*ڊ�6�<�;�
��}�JϽ�&����l��Z1�����=�&���$�>�F�������]ǑN��X���
�
�6�<�9��(߁�	������^	�����0�&�u�x�w�}����8����]��h^�����1�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���K����lT��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��_��\ʡ�0�u�u�u�w�}�W���	�֓�P��Y��*ڊ�%�#�1�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����lV��T�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�e��)�������F��h �����'�
�=�0��<����&����9��P1�E��_�u�u�x�'�m�6�������lW��G1��ʴ�&�2�u�'�4�.�Y��s���C9��v�����0�d�4�
�;���������PF��G�����4�
�0�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�d�|�u�?�3�}���Y���F�G1��4���:�&�0�d�6�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N������!�:�&�2�l���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W���&����\��R1�I���9�;�1�
�2�0�4�������\��X��*���
�b�c�_�w�}�Z���&ù��G��D1��G���
�9�u�&�>�3�������KǻN��*ڊ�6�<�;�
����������Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�d�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�e�t�^Ϫ���ƹF�N��U���
�
�6�<�9��(݁�	����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�
�4�4����&����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����lV��T�����
�u�h�6��2��������@��R
�����9�&�d�'�0�l�E��s���K��h^�����;�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�e��)�����Փ�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!�e�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���F��R ��U���u�u�u�u�'�m�6�������lU��G1����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����8����]��h]�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN������!�:�&�2�i�K�������V9��E�����1�1�:�!�8��(݁�����P��=N��U���%�e��!�8�.��������WF��D��U���6�&�{�x�]�}�W���&����\��R1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K����^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h\�\���=�;�_�u�w�}�W���Y����r��X �����4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��v�����0�a�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
��>����&����[��[1�����0�8��&�6�8�4�������lU��R	��B��_�u�u�x�w��(�������V9��V�����&�<�;�%�8�8����T�����h/�����
�
�
�%�!�9��������\������}�%�6�y�6�����
����g9��\�����d�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��G���8�g�|�|�#�8�W���Y���F���*���<�;�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���
�6�<�;���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�I����Z	��h��U��6�
�:�0�#�/�(�������p	��E�����'�2�d�f�l�W�W���TӖ��l'��^��*���
�%�#�1�6�.��������@H�d��Uʥ�e��!�:�$�8�A���&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�g�3�8�e�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��F���Y����l�N��U���u�%�e��#�2����O����E
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�%�g�����
����l��A��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��1�����&�0�b�i�w�1����&����l%��T�����!�:�
�
��8�(��H��ƹF�N��E���!�:�&�0�`�<�(���Y����T��E�����x�_�u�u����������9��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�o�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O����ߊu�u�u�u�w�}�(߁�����@9�� 1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&ù��G��D1��B���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�
�6�<�9��(���DӅ��]	��h�����&�4�0��9�/����O����lW��UװU���x�u�
�
�4�4����&˹��l�������%�:�0�&�w�p�W���	�֓�P��Y��*Ҋ�%�#�1�4�$�:�(�������A	��D�����y�4�
�<��.����&����l ��h\����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���|�!�0�u�w�}�W���Y����lV��T�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��h^�����;�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�m�6�������l_�
N��*���0�!�'�
�6�>��������_9�� 1����`�n�_�u�w�p����8����]��hW�����1�4�&�2�w�/����W���F�G1��4���:�&�0�l�6�����
����l��TN����0�&�4�
�2�}��������B9��h��G���8�g�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�}����s���F�N������!�:�&�2�d���������T�����2�6�d�_�w�}�W������F�N��U���%�e��!�8�.��������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��h=�����!�
�
�
�'�+����&����R��P �����&�{�x�_�w�}�(���*����Z��h��*���#�1�<�
�>���������PF��G�����%�d�
�0�'�4����&ù��l��N��Dڊ�0�%�<�!���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�d�
�2�-����&����R��[
��U���;�_�u�u�w�}�W���&�֓�V��^ ��*���
�%�#�1�>�����DӖ��9��C�����0�e�4�
�;�f�W���Y����_��=N��U���u�u�u�
�g���������lV��G1�����
�<�u�h�'�l�(���	����@9��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����l5��G�����
�
�;�&�0�<����Y����V��C�U���%�d�
�0�'�4����&ù��l��h�����%�:�u�u�%�>����&�֓�V��^ ��*���y�%�d�
�2�-����&����C��N��Dڊ�0�%�<�!���(������F�U�����u�u�u�<�w�u��������\��h_��U���e��!�:�9�.��������WO�C��U���u�u�u�u�w�-�F߁�����]��R1�����<�u�h�%�f���������V9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�V��R�����
�
�
�;�$�:�K���&�֓�V��^ ��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����l/��B�����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�d��3�����֓�C9��S1��*���
�&�<�;�'�2�W�������@N��_�����&�0�e�4��1�[Ϯ�H¹��C��h��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�W��Y�����e�4�
�9�~�}����s���F�N����
�;� �&�2�m��������l��R����
�;� �&�2�m������ƹF�N�����_�u�u�u�w�}�W���H����F��R1�����9�
�;�&�0�a�W���H����F��R1�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�W��Y�����e�<�
�<�w�.����	����@�CךU���
�d��%�#��(߁�����l��^	�����u�u�'�6�$�u�(���0����@9��B��*����%�!�
������Y����l/��B�����4�
�9�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����l/��B�����4�
�9�|�w�5��ԜY���F�N��Dۊ�;� �&�0�g�4�(���Y����lW��~ �����
�n�u�u�w�}����Y���F�N��U���d��%�!���(���
���F��_�����&�0�e�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����1�����
�
�
�%�!�9�����ƭ�@�������{�x�_�u�w��F���	����V9��V�����;�&�2�4�$�:�(�������A	��D��*����%�!�
�������Ƽ�W��Y�����d�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h_��<���!�
�
�
�'�+��������9F�N��U���u�
�d��'�)�(���&����_��Y1����u�
�d��'�)�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��9��G��*���
�%�#�1�>�����DӖ��9��G��*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h_��<���!�
�
�
�9�.�Ͽ�
����C��R��U���u�u�%�d��3�����ד�]9��P1�����
�'�6�o�'�2����	����z��C��*���%�d�
�;�"�.����	������1�����
�
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������1�����
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�d��%�#��(ށ�����Z�G1�*��� �&�0�d�]�}�W���Y����l�N��U���u�%�d�
�9�(����H����@��S��*����%�!�
������s���F�R ����_�u�u�;�w�/����B��ƹF�N��Dۊ�;� �&�0�e�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�H¹��C��h��*���#�1�<�
�>���������PF��G�����%�d�
�;�"�.��������WJ��h_��<���!�
�
�
�'�+������ƹF��R	�����u�u�u�3��<�(���
����T��N����
�;� �&�2�o�������G��d��U���u�u�u�%�f�����
����l��A�����<�u�h�%�f�����
����l��A�����u�u�u�9�2�W�W���Y���F��_�����&�0�g�4��1�(���
���F��_�����&�0�g�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C���
�;� �&�2�o�����ƭ�@�������{�x�_�u�w��F���	����V9��^ �����&�<�;�%�8�}�W�������C9��h'�� ���0�g�u�
�f�����&����C��N��Dۊ�;� �&�0�e�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��Dۊ�;� �&�0�e�<�(���P�Ƹ�V�N��U���u�u�%�d��3�����ԓ�]9��PN�U���d��%�!���L���Y�����RNךU���u�u�u�u��l�>�������9��h��U��%�d�
�;�"�.����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�d��%�#��(܁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�W��Y�����f�4�
�9��3��������]9��X��U���6�&�}�
�f�����&����R��[
���
�;� �&�2�n��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�d��'�)�(���&����_����ߊu�u�u�u�w�}�(���0����@9��1��*���
�;�&�2�k�}�(���0����@9��1��*���n�u�u�u�w�8����Y���F�N��*����%�!�
����������@��S��*����%�!�
����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�d��'�)�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�H¹��C��h��*���&�2�4�&�0�����CӖ��P����D���%�!�
�
�{�-�Fށ�����l��h�����
�d��%�#��(܁�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�d��%�#��(܁�	����O��_�����u�u�u�u�w��F���	����V9��^ �����h�%�d�
�9�(����J���F�N�����u�u�u�u�w�}���&����G��h]�����2�i�u�
�f�����&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�d��3�����ғ�C9��S1��*���u�&�<�;�'�2����Y��ƹF��h_��<���!�
�
�
�'�+����&����R��P �����o�%�:�0�$�-�Fށ�����l��h�����u�
�d��'�)�(���&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�f�����
����l��A��\ʡ�0�u�u�u�w�}�W���	����z��C��*ފ�%�#�1�<��4�W��	����z��C��*ފ�%�#�1�_�w�}�W������F�N��U���%�d�
�;�"�.��������W9��h��U��%�d�
�;�"�.��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�f�����
����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�W��Y�����a�<�
�<��.����	����	F��X��¥�d�
�;� �$�8�C���&�ד�]��D1��A���0�y�%�d��3�����ғ�C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�d��3�����ғ�C9��SG�����u�u�u�u�w�}�WϮ�H¹��C��h��*���&�2�i�u��l�>�������]ǻN��U���9�0�_�u�w�}�W���Y����l/��B�����<�
�<�u�j�-�Fށ�����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��F���	����V9��V�����;�&�2�4�$�:�W�������K��N����
�;� �&�2�h��������l��h�����%�:�u�u�%�>����&�ד�]��D1��@���
�9�y�%�f�����
����l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(���0����@9��1��*���|�u�=�;�]�}�W���Y���C9��h'�� ���0�`�4�
�;��������C9��h'�� ���0�`�4�
�;�f�W���Y����_��=N��U���u�u�u�
�f�����&����R��[
�����2�i�u�
�f�����&����R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(���0����@9��1��*���u�&�<�;�'�2����Y��ƹF��h_��<���!�
�
�
�9�.����
����C��T�����&�}�
�d��-����&����lW��~ �����
�
�'�2�w��F���	����V9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��F���	����V9��V�����u�=�;�_�w�}�W���Y�Ƽ�W��Y�����`�<�
�<�w�`���&����G��h[�U���u�u�0�&�w�}�W���Y�����1�����
�
�
�;�$�:�K���&�ד�]��D1��@���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�H¹��C��h��*���#�1�<�
�>�}����Ӗ��P��N����u�
�d��'�)�(���&����_��Y1�����&�2�
�'�4�g��������lW��~ �����
�
�%�#�3�}�(���0����@9��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	����z��C��*܊�%�#�1�|�#�8�W���Y���F���D���%�!�
�
��-��������TF���D���%�!�
�
��-����s���F�R��U���u�u�u�u�w�-�Fށ�����l��h�����<�
�<�u�j�-�Fށ�����l��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	����z��C��*܊�;�&�2�4�$�:�W�������K��N����
�;� �&�2�k��������@��h����%�:�0�&�'�l�(�������lP�G1�*��� �&�0�c�'�8�[Ϯ�H¹��C��h��*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�H¹��C��h��*���#�1�|�!�2�}�W���Y���F��h_��<���!�
�
�
�9�.���Y����l/��B����_�u�u�u�w�1��ԜY���F�N��Dۊ�;� �&�0�a�4�(���Y����lW��~ �����
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���&����G��D1��E��u��-� �.�(�(ց�����P��=N��U���%�f��!�"�.��������WF��D��U���6�&�{�x�]�}�W���&����F��R1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K����^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h\�\���=�;�_�u�w�}�W���Y����|��B�����4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��x�� ���0�e�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
��(����&����[��E�� ��b�%�n�u�w�-�D�������l��N�U�������8�)����N����l��h_�L�ߠu�u�x�u����������V��G1��ʴ�&�2�u�'�4�.�Y��s���C9��x�� ���0�d�
�%�!�9��������\������}�%�6�y�6�����
����g9��\�����d�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��G���8�g�|�|�#�8�W���Y���F���*���%�!�
�
�g�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�f��!� �$�8�F߁�	����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lU��B�����
�
�%�#�3�<����Y����V��C�U���%�f��!�"�.��������W9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�g�3�:�o�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�g��.�(��P�Ƹ�V�N��U���u�u�%�f��)�����ד�C9��SN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�'�n�8�������lW��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�G1��:��� �&�0�g�k�}��������l��=d��U���u�
�
� �'�)�(���&����_��D��ʥ�:�0�&�u�z�}�WϮ�J����C��h��*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ԓ�@��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӖ��l)��G��*���
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����h!�����
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�%�d�����
����Z�Q=��&����!�l�'�0�l�B��s���K��h]�� ���!�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�f��)�����Փ�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!�e�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���F��R ��U���u�u�u�u�'�n�8�������lU��G1����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����6����G��h]�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN������!� �&�2�i�K���*����w��C1�����d�c�n�_�w�}�ZϮ�J����C��h��*���#�1�4�&�0�}����
���l�N��F���!� �&�0�c�<�(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�g�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�f�t�W������F�N��Uʥ�f��!� �$�8�C���&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�%�f��#�(����M����E
��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�Ƽ� 9��C�����`�i�u�0��o�L�ԜY�����h!�����
�
�
�%�!�9�����Ƽ�\��D@��X���u�%�f��#�(����L����E
��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�g�1�0�E���Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�e�����H���G��d��U���u�u�u�%�d�����
����l��A��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�-�D�������l��h�����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N��F���!� �&�0�a�a�W���&����9l�N�U���
� �%�!���(�������@��YN�����&�u�x�u�w�-�D�������l��h�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���K����^9��G�����u�u�u�u�w�}�WϮ�J����C��h��*���#�1�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӖ��l)��G��*���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�f��#�(����N���U5��v*��:���g�
�
�0��k�O�ԶY���F��1�����&�0�b�4��1�W�������A	��D�X�ߊu�u�
�
�"�-����&Ĺ��l��h�����%�:�u�u�%�>����	������D�����
��&�g��.�(��s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�o����K�����YNךU���u�u�u�u����������9��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}�(܁�����@9�� 1��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN��*ي� �%�!�
��}�Jϸ�&����J)��h=�����!�d�
�
�2��A��s���K�G1��:��� �&�0�m�6�����
������T��[���_�u�u�
��(����&����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�����H���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�E�������O��_�����u�u�u�u�w��(���	����V9��V�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����F��R1�����9�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=N��U���
� �%�!���W������W��R��!���0�=�&���.��������]ǑN��X���
�
� �%�#��(ց�	������^	�����0�&�u�x�w�}����6����G��hW�����1�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���K����lT��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��_��\ʡ�0�u�u�u�w�}�W���	�Փ�F��C��*ӊ�%�#�1�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����lU��B�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�i�:�������G��h��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�4�"�1��������9��h��*���&�2�4�&�0�����CӖ��P����*��� �9�:�!�8��(߁�	����F��1������;�'�9�2�m��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�4�"�1��������9��h��\���=�;�_�u�w�}�W���Y����~��V�����9�0�e�4��1�(���
���F��1������;�'�9�2�m������ƹF�N�����_�u�u�u�w�}�W���&����R
��Y�����e�4�
�9��3����E�Ƽ�9��Y��6���'�9�0�e�6���������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�a��;�4��3�����֓�]9��PN�����u�'�6�&�y�p�}���Y����~��V�����9�0�e�<��4�(�������A	��N�����&�%�a��9�<�4�������lV�G1��8���4��;�'�;�8�G�������lR��V �����!�:�
�
��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*��� �9�:�!�8��(߁�	����O��_�����u�u�u�u�w��(�������]��[1��E���
�<�u�h�'�i�:�������G��h��N���u�u�u�0�$�}�W���Y���F��hZ�����9�:�!�:���(���
���F��1������;�'�9�2�m����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ފ�4� �9�:�#�2�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��z�����;�'�9�0�f�<�(���&����Z��D�����:�u�u�'�4�.�_���&����R
��Y�����d�4�
�9�{�-�C�������\��X��*ۊ�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��z�����;�'�9�0�f�<�(���P�Ƹ�V�N��U���u�u�%�a��3��������l��h�����<�
�<�u�j�-�C�������\��X��*ۊ�%�#�1�_�w�}�W������F�N��U���%�a��;�6���������l��A�����<�u�h�%�c�����:����\
��h_�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l+��B�����:�
�
�
�9�.�Ͽ�
����C��R��U���u�u�%�a��3��������l��h�����4�&�2�
�%�>�MϮ�������h#�� ���:�!�:�
��q����4����_%��C��*���
�'�2�u����������A	��R1�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R
��Y�����d�4�
�9�~�}����s���F�N������;�4��9�/����H����@��S��*ފ�4� �9�:�#�2�(���B���F����ߊu�u�u�u�w�}�(ہ�����p	��E�����<�
�<�u�j�-�C�������\��X��*ۊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ǹ��]��t�����0�g�4�
�;�����Ӈ��Z��G�����u�x�u�u�'�i�:�������G��h��*���#�1�<�
�>���������PF��G�����%�a��;�6���������l��A��U���
�4� �9�8�)����&����l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�i�:�������G��h��*���#�1�|�!�2�}�W���Y���F��hZ�����9�:�!�:���(�������]9��PN�U���
�4� �9�8�)����&����l��d��U���u�0�&�u�w�}�W���Y����lR��V �����!�:�
�
��-��������TF���*��� �9�:�!�8��(݁�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��<��������_9��1��*���u�&�<�;�'�2����Y��ƹF��hZ�����9�:�!�:���(���
����@��Y1�����u�'�6�&���(�������]��[1��G���
�
�4� �;�2����&����C��N��A���;�4��;�%�1��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�a��;�6���������l��A��\ʡ�0�u�u�u�w�}�W���	�ғ�R��[-�����
�
�
�;�$�:�K���&ǹ��]��t�����0�g�_�u�w�}�W������F�N��Uʥ�a��;�4��3�����ԓ�]9��PN�U���
�4� �9�8�)����&����V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�a��9�<�4�������lU��G1�����
�<�u�&�>�3�������KǻN��*ފ�4� �9�:�#�2�(���&����_��Y1�����&�2�
�'�4�g��������lR��V �����!�:�
�
��-����Y����~��V�����9�0�f�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ފ�4� �9�:�#�2�(���&����_����ߊu�u�u�u�w�}�(ہ�����p	��E�����4�
�9�
�9�.���Y����~��V�����9�0�f�4��1�L���Y�����RNךU���u�u�u�u����������A	��R1�����9�
�;�&�0�a�W���&����R
��Y�����f�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��8���4��;�'�;�8�D���&����R��P �����&�{�x�_�w�}�(ہ�����p	��E�����<�
�<�
�$�4��������C��R������;�4��9�/����J�Ƽ�9��Y��6���'�9�0�f�'�8�[Ϯ�M����F��X �����
�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lR��V �����!�:�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�(��������V9��^ �����h�%�a��9�<�4�������lU��N��U���0�&�u�u�w�}�W���YӖ��l+��B�����:�
�
�
�9�.���Y����~��V�����9�0�f�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h#�� ���:�!�:�
����������@��V�����'�6�&�{�z�W�W���&ǹ��]��t�����0�a�4�
�;���������Z��G��U���'�6�&�}����������A	��R1�����9�y�%�a��3��������l��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ǹ��]��t�����0�a�4�
�;�t�W������F�N��Uʥ�a��;�4��3�����ғ�C9��S1��*���u�h�%�a��3��������l��h�����_�u�u�u�w�1��ԜY���F�N��A���;�4��;�%�1��������W9��h��U��%�a��;�6���������l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����4����_%��C��*���
�;�&�2�6�.��������@H�d��Uʥ�a��;�4��3�����ғ�]9��P1�����
�'�6�o�'�2����	�ғ�R��[-�����
�
�y�%�c�����:����\
��hZ�����u�
�
�4�"�1��������9��h��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u����������A	��R1�����9�|�u�=�9�W�W���Y���F��1������;�'�9�2�i���������h#�� ���:�!�:�
��f�W���Y����_��=N��U���u�u�u�
��<��������_9��1��*���u�h�%�a��3��������l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������]��[1��@���
�9�
�;�$�:�����Ƽ�\��D@��X���u�%�a��9�<�4�������lS��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��A���;�4��;�%�1��������WJ��hZ�����9�:�!�:���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�a��9�<�4�������lS��G1�����!�0�u�u�w�}�W���YӖ��l+��B�����:�
�
�
�'�+����&����[��hZ�����9�:�!�:���(�������F�N�����u�u�u�u�w�}�WϮ�M����F��X �����
�
�%�#�3�4�(���Y����lR��V �����!�:�
�
��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�4� �;�2����&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l+��B�����:�
�
�
�9�.����
����C��T�����&�}�
�
�6�(��������V9����*��� �9�:�!�8��(ځ����C9��z�����;�'�9�0�b�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��A���;�4��;�%�1��������WO�C��U���u�u�u�u�w�-�C�������\��X��*ߊ�;�&�2�i�w��(�������]��[1��@�ߊu�u�u�u�;�8�}���Y���F�G1��8���4��;�'�;�8�B���&����[��hZ�����9�:�!�:���(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C�����;�4��9�/����O����E
��^ �����&�<�;�%�8�8����T�����h#�� ���:�!�:�
����������@��V�����'�6�o�%�8�8�Ǯ�M����F��X �����
�
�%�#�3�}�(ہ�����p	��E�����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h#�� ���:�!�:�
����������[��=N��U���u�u�u�
��<��������_9��1��*���
�;�&�2�k�}�(ہ�����p	��E�����4�
�9�n�w�}�W�������9F�N��U���u�
�
�4�"�1��������9��h��*���&�2�i�u����������A	��R1�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Y��6���'�9�0�c�>�����
������T��[���_�u�u�
��<��������_9��1��*���
�&�<�;�'�2�W�������@N��1������;�'�9�2�k�W���&����R
��Y�����c�%�0�y�'�i�:�������G��h��*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�M����F��X �����
�
�%�#�3�t����Y���F�N��U���
�4� �9�8�)����&Ź��l��R������;�4��9�/����O���F�N�����u�u�u�u�w�}����4����_%��C��*���
�;�&�2�k�}�(ہ�����p	��E�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ғ�R��[-�����
�
�
�%�!�9�����ƭ�@�������{�x�_�u�w��(�������]��[1��B���
�9�
�;�$�:��������\������}�
�
�4�"�1��������9��h��Yʥ�a��;�4��3�����ѓ�C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(�������]��[1��B���
�9�|�u�?�3�}���Y���F�G1��8���4��;�'�;�8�@���&����Z��^	��Hʥ�a��;�4��3�����ѓ�C9��SUךU���u�u�9�0�]�}�W���Y���C9��z�����;�'�9�0�`�<�(���&����Z�
N��A���;�4��;�%�1��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�c�����:����\
��hY�����2�4�&�2�w�/����W���F�G1��8���4��;�'�;�8�@���&����R��P �����o�%�:�0�$�-�C�������\��X��*���%�a��;�6���������l��PB��*ފ�4� �9�:�#�2�(���&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�4�"�1��������9��h��\���=�;�_�u�w�}�W���Y����~��V�����9�0�b�<��4�W��	�ғ�R��[-�����
�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�4� �;�2����&����Z��^	��Hʥ�a��;�4��3�����ѓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����e�4�
�9��3��������]9��X��U���6�&�}�
��<����&ù��l��N��@���;�0�0�e�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&ù��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*ڊ�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�m��������@��h����%�:�0�&�'�h�%�������F��1�����0�e�%�0�{�-�B�������lV��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������֓�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����d�4�
�9��3��������]9��X��U���6�&�}�
��<����&¹��l��N��@���;�0�0�d�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&¹��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*ۊ�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�l��������@��h����%�:�0�&�'�h�%�������F��1�����0�d�%�0�{�-�B�������lW��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������ד�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����g�4�
�9��3��������]9��X��U���6�&�}�
��<����&����l��N��@���;�0�0�g�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&����l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*؊�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�o��������@��h����%�:�0�&�'�h�%�������F��1�����0�g�%�0�{�-�B�������lT��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������ԓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����f�4�
�9��3��������]9��X��U���6�&�}�
��<����&����l��N��@���;�0�0�f�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&����l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*ي�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�n��������@��h����%�:�0�&�'�h�%�������F��1�����0�f�%�0�{�-�B�������lU��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������Փ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����a�4�
�9��3��������]9��X��U���6�&�}�
��<����&ǹ��l��N��@���;�0�0�a�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&ǹ��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*ފ�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�i��������@��h����%�:�0�&�'�h�%�������F��1�����0�a�%�0�{�-�B�������lR��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������ғ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����`�4�
�9��3��������]9��X��U���6�&�}�
��<����&ƹ��l��N��@���;�0�0�`�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&ƹ��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*ߊ�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�h��������@��h����%�:�0�&�'�h�%�������F��1�����0�`�%�0�{�-�B�������lS��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������ӓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����c�4�
�9��3��������]9��X��U���6�&�}�
��<����&Ź��l��N��@���;�0�0�c�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&Ź��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*܊�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�k��������@��h����%�:�0�&�'�h�%�������F��1�����0�c�%�0�{�-�B�������lP��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������Г�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����b�4�
�9��3��������]9��X��U���6�&�}�
��<����&Ĺ��l��N��@���;�0�0�b�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&Ĺ��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*݊�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�j��������@��h����%�:�0�&�'�h�%�������F��1�����0�b�%�0�{�-�B�������lQ��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������ѓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����m�4�
�9��3��������]9��X��U���6�&�}�
��<����&˹��l��N��@���;�0�0�m�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&˹��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*Ҋ�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�e��������@��h����%�:�0�&�'�h�%�������F��1�����0�m�%�0�{�-�B�������l^��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������ޓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�:�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e�����l�4�
�9��3��������]9��X��U���6�&�}�
��<����&ʹ��l��N��@���;�0�0�l�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�2�
����������[��=N��U���u�u�u�
��<����&ʹ��l��h�����i�u�
�
�6�:�(���&����_��N��U���0�&�u�u�w�}�W���YӖ��l4��P��*ӊ�%�#�1�<��4�W��	�ӓ�R��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lS��V ��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�d��������@��h����%�:�0�&�'�h�%�������F��1�����0�l�%�0�{�-�B�������l_��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�%�������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�R��h��*���&�2�i�u������&����9F�N��U���0�_�u�u�w�}�W���&ƹ��]��R1�����<�u�h�%�b������ߓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�<����
����l��A�����<�u�&�<�9�-����
���9F���*���4�0�0�&�2�m��������l��h�����%�:�u�u�%�>����&Ź��A��C��*���
�%�#�1�w��(�������A��h^�����1�%�0�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����c��Z�����
�
�%�#�3�t����Y���F�N��U���
�4�4�0�2�.��������W9��h��U��%�c��'�:�)����&ù��l��d��U���u�0�&�u�w�}�W���Y����lP��V�����&�0�e�4��1�(���
���F��1�����!�'�
�
��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�4�4�2�8����I����@��V�����'�6�&�{�z�W�W���&Ź��A��C��*���
�;�&�2�6�.���������T��]���
�4�4�0�2�.���Y����c��Z�����
�
�'�2�w��(�������A��h^�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����)����V��D1��E���
�9�|�u�?�3�}���Y���F�G1��%���8�!�'�
���������C9��g�����'�
�
�n�w�}�W�������9F�N��U���u�
�
�4�6�8�����֓�]9��PN�U���
�4�4�0�2�.����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�4�4�2�8����H����E
��^ �����&�<�;�%�8�8����T�����h>�����0�&�0�d�6���������l��^	�����u�u�'�6�$�u�(ف�����G��h��*���#�1�u�
��<��������lW��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����^��E��*ۊ�%�#�1�|�#�8�W���Y���F���*���4�0�0�&�2�l��������l��R������'�8�!�%��(ށ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�Г�R��R�����d�4�
�9��3����E�Ƽ�9��E�����
�
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*܊�4�4�0�0�$�8�F���&����R��P �����&�{�x�_�w�}�(ف�����G��h��*���&�2�4�&�0�����CӖ��P����*���4�0�0�&�2�l�W���&����^��E��*ۊ�'�2�u�
��<��������lW��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�k�'�������@9��1��*���|�u�=�;�]�}�W���Y���C9��g�����'�
�
�
�9�.���Y����c��Z�����
�n�u�u�w�}����Y���F�N��U���
�4�4�0�2�.��������TF���*���4�0�0�&�2�l����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lV��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�e�<�
�>���������PF��G�����%�b��<�$�8�G���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�G���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�m����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lW��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�d�<�
�>���������PF��G�����%�b��<�$�8�F���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�F���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�l����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lT��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�g�<�
�>���������PF��G�����%�b��<�$�8�E���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�E���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�o����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lU��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�f�<�
�>���������PF��G�����%�b��<�$�8�D���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�D���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�n����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lR��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�a�<�
�>���������PF��G�����%�b��<�$�8�C���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�C���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�i����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lS��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�`�<�
�>���������PF��G�����%�b��<�$�8�B���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�B���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�h����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lP��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�c�<�
�>���������PF��G�����%�b��<�$�8�A���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�A���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�k����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9�� 1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������lQ��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�b�<�
�>���������PF��G�����%�b��<�$�8�@���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�@���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�j����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������l^��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�m�<�
�>���������PF��G�����%�b��<�$�8�O���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�O���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�e����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�;�&�2�6�.���������T��]���
�4�;�
�������Ƽ�9��^ �����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h)�����
�
�%�#�3�t����Y���F�N��U���
�4�;�
����������@��S��*݊�4�;�
�
��-����s���F�R��U���u�u�u�u�w�-�@�������l_��G1�����
�<�u�h�'�j�0���
����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����>����l��h�����4�&�2�u�%�>���T���F�� 1�����0�l�<�
�>���������PF��G�����%�b��<�$�8�N���&Ĺ��Z��R1�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��<�$�8�N���&����F��R ��U���u�u�u�u�'�j�0���
����l��D��I���
�
�4�;���L���Y�����RNךU���u�u�u�u������&����Z��^	��Hʥ�b��<�&�2�d����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ӊ�<�;�9�
����������@��V�����'�6�&�{�z�W�W���&ʹ��T��D1��E���
�9�
�;�$�:��������\������}�
�
�<�9�1�(���&����_�G1��&���4�&�0�e�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�<�;�9���(��������YNךU���u�u�u�u����������9��h��*���&�2�i�u����������9��h��N���u�u�u�0�$�}�W���Y���F��hW�����9�
�
�
�'�+����&����[��hW�����9�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�<�;�9���(���
����@��YN�����&�u�x�u�w�-�N�������l��h�����4�&�2�
�%�>�MϮ�������h=�����
�
�y�%�n�����
����l��PB��*ӊ�<�;�9�
���������F��P��U���u�u�<�u��-��������Z��S��*ӊ�<�;�9�
����������[��=N��U���u�u�u�
��4����&����Z��^	��Hʥ�l��2�4�$�8�G�ԜY���F��D��U���u�u�u�u�'�d�$�������lV��Y1����u�
�
�<�9�1�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�l��2�6�.��������W9��h��U���<�;�%�:�2�.�W��Y����l_��^	�����
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�n�����
����l��A��U���
�<�;�9���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�l��0�<����H����E
��N�����u�u�u�u�w�}����*����_��h_�����1�<�
�<�w�`����*����_��h_�����1�_�u�u�w�}����s���F�N������2�4�&�2�l��������l��R������2�4�&�2�l��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�l��0�<����H����@��V�����'�6�&�{�z�W�W���&ʹ��T��D1��D���
�<�
�&�>�3����Y�Ƽ�\��DF��L���2�4�&�0�f�}�(ց�����@9��1�����%�l��2�6�.��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�l��2�6�.��������WO�C��U���u�u�u�u�w�-�N�������l��h�����i�u�
�
�>�3����&��ƹF�N�����_�u�u�u�w�}�W���&����R
��R1�����<�u�h�%�n�����
����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�
�0� �#�e�(���A�ד� F�F��*���&�
�#�e�g�{����/����^��GZ����u�
�0� �#�e�(���@�ߓ�F�F��#���
�
� �b�f�-�_������\F��N�����b�
�
� �n�l����s���C9��D��*���3�
�e�d�'�}�J���	����@��A_��E��9�6��g��(�N���	����F�G1�����
�e�3�
�f�d����D�μ�e��hY�����b�
�d�f�w�2����J�����hY��ۊ� �d�d�
�d�f�W���	����F
��_�� ��m�
�`�i�w�-�!���&�ד�F9��_��D��u�:�;�:�d�t�QϪ�	����Z9��h_�E���|�_�u�u��8����
����U��h�I���4�
�:�&��+�G��_ӊ��l0��1��*��a�%�|�_�w�}�(���K����U�� _��D��u�
�d��'�)�(���&����Z��N�����9�
�d�3��o�F���Y����`9��b,�� ���
�0�
�b�a�W�W���&����l��B1�D���u�h�%�d��3�����֓�]9��PUךU���0�
�
�
��i�(�������G9��h_�A���u�h�_�u�w�}�W�������l
��1�Eʢ�0�u�!�%�>�4�ށ�I����T��h�E���u�d�|�0�$�}�W���Y����C9��Y����
�e�n�u�w�/��������
9��D�����3�
�e�`�'�}�J�ԜY���F��h�����#�`�`�e� �8�WǪ�	����l��Q��Lߊ�g�e�u�u�f�t����Y���F������!�9�d�
�g�f�W�������l��h�����6�&�
� �o�h����D���F�N��*���&�
�#�`�b�m� ���Yے��l��h��L���
�e�
�g�g�}�W��PӃ��VFǻN��U���%�6�;�!�;�l�(��B�����h��*���3�
�g�e�'�}�J�ԜY���F��h�����#�`�a�e�w�5��������Z9��hZ�����g�a�%�}�~�`�P���Y����l�N��Uʴ�
�:�&�
�!�h�C��B�����h��*���3�
�e�d�'�}�J�ԜY���F��h�����#�`�a�e�w�5��������Z9��h��L���%�}�|�h�p�z�W������F�N��*���&�
�#�`�c�m�L���YӔ��l��h�� ��d�%�u�h�]�}�W���Y����\��h��@��e�u�=�;��0�(���&����l ��^�����|�h�r�r�w�1��ԜY���F��h�����#�`�a�e�l�}�Wϭ�����9��h��D��
�g�i�u�#�-����ƹ��l_��h����4�
�:�&��+�(���s���@��C��*���3�
�f�e�'�}�J�������Z9��h��D���
�g�-�'�6�����&����O��N�����!�%�
�
�"�e�F���Y���G��^1�����
�l�
�g�/�/��������_��G�U���&�9�!�%��i����I�ѓ�F�F����b�<�<�<��(�F��&����]��R�����<�
� �d�d��E��Y����V
��Z��ߊ� �d�e�
�e�a�WǪ�	����l��h�����g�m�%�u�9�}�����ד�9��h_�E���|�_�u�u�2���������R��G\��H���8�
�f�
���(���A�ߓ�F��SN�����%�
�
� �o�l����s���@��C��*���3�
�d�`�'�}�J���[ӑ��]F��d1�� ���;� �
�e�>������ד�F9��]��F��4�
�:�&��+�B��I����_��^�����u�0�
�8�a�4�(���H����CT�
N��Wʢ�0�u�3�
���E����ѓ�]9��c��*���d�d�
�f�j�<�(���
����S��^�U���0�w�w�_�w�}�����Г�l ��Z�����h�w�w�"�2�}����4����])��h\�����%�,�0�3��h�(��DӇ��P	��C1��Dߊ�a�e�u�9�2��U�ԜY�ƿ�_9��GY��D���
�d�d�%�w�`�U������� ��O#��!ػ� �
�e�<��-����H����V��h�Hʴ�
�:�&�
�!�h�C��Y����D��d��Uʦ�9�!�%�
�e�;�(��I����[�L�����}��-� ��3����&����C2��R1��*��g�%�u�u�'�>��������V�������w�_�u�u�2���������
S��G\��H���w�"�0�u�1��:���K����lT��^ �����0�3�
�`��n�JϿ�&����G9��[��E���0�&�u�e�l�}�Wϭ�����9��h��D��
�g�i�u�$�1����&�ԓ�F9��[��Gʺ�u�0�
�8�`�4�(���H����CT�=N��U���
�8�m�<��(�F��&���F��R�����<�
� �d�g��Eϱ�Y����G��h�����a�e�%�|�]�}�W���&����l��B1�B���u�h�}�0��0�A�������9�������!�%�
�
�"�d�F���P���F��[1�����
� �d�g��n�K���Y���F��R��*���b�3�
�e�f�-�W����θ�C9��^1��*���l�l�%�}�~�`�P���Y����l�N��Uʴ�
�:�&�
�!�h�C��s���@��C��ߊ� �d�l�
�d�a�W���Y�����h��*���3�
�g�e�'�}����Q����Z9��^_�� ��`�
�g�e�w�}�F�������9F�N��U���6�;�!�9�f��G��Y����V
��Z��*���m�f�%�u�j�W�W���Y�ƾ�G9��^1�����d�
�f�"�2�}��������l �� W�����|�h�r�r�w�1��ԜY���F��h�����#�`�a�e�]�}�W���&����ZW��B1�Bۊ�g�i�u�d�w�5�������� ��O#��!ػ� �
�e�<��%�(���&����S��G\��Iʦ�2�0�}�%�4�3����H˹��F��D��E��u�u�!�%�f�m����&����CT�
N��Wʢ�0�u�&�2�2�u�$���,����|��^�����%��d�3��k�(��Y�ƿ�T�������!�9�d�
�~�}����[����F�C��D���3�
�e�
�f�a�W���������C1�*���0�%��d�1��Aց�K���W��X����n�u�u�!�'�l�C���&����l��S��&��� ��;� ��m�������� 9��h_�L���}�u�u�u�8�3���B�����h_�*���d�c�
�d�k�}�$���,����|�� 1��*���
�
�
� �f�o�(��A�����Y��E��u�u�!�%�f�n����&����l��S��D���=�;�}�<�9�9����4����])��hY�����%��d�3��n�O���P����Z��SF��*���&�
�#�m�f�t����Y���9F���*��
�
�
�d�1��E���	���D�������:�
�
�g�1��E���	���R��X ��*���
��u�9�2��U�ԜY�Ƹ�C9�� 1�����
� �d�e��o�K���H�ƻ�V�[��#��
� �l�`�'�}�W�������l
��h(��U���0�w�w�_�w�}����JĹ��Z9��Q��Dӊ�g�i�u�d�w�5��������U��[��A��4�
�:�&��+�(���Y����D��d��Uʡ�%�c�
� �n�l����D���F�N��*���&�
�#�
��*��������l ��Y�����|�h�r�r�w�1��ԜY���F��h�����#�
�n�u�w�)���&����_��G]��H�ߊu�u�u�u�'�>�����ޓ�uF��R �����<�
� �d�a��E��Y���O��[�����u�u�u�%�4�3����A����F�C��Cߊ� �d�c�
�d�a�W���Y�����T�����m��u�=�9�u����J����U��h�E���u�d�|�0�$�}�W���Y����C9��Y�����e�_�u�u�:��C���&����W��G]��H���8�
�f�3��l�D���Y�Ƽ�T��h_��D���
�e�f�%�~�W�W�������l��B1�D���u�h�}�8��l����H����@��h^�E���<�3�
�l��n�L���YӒ��l^��Q��Dي�f�i�u�u�w�}�WϪ�	����U��_��Fʢ�0�u�!�%�1��O؁�K���F�G�����_�u�u�u�w�0�(��&����_��UךU���8�
�g�3��m�@���Y���G��^\�� ��c�
�g�:�w�0�(��&�ד�F9�� _��G��u�u�!�%�o����I����Z�=N��U���u�8�
�a�1��G���	�ƻ�V�C��M؊� �d�b�
�e�m�W���H����_��=N��U���u�8�
�e��(�F��&����F�C��Mފ� �d�a�
�e�a�WǪ�	����U��]�����'�!�%�d�d�4����J�֓�O��N�����m�
� �d�`��D��Y���F���*���3�
�f�e�'�}����Q����R��B1�A܊�g�e�u�u�f�t����Y���F���*��
� �d�c��l�}���Y����Q��h��D��
�f�i�u�#�-�Oځ�����9��H��*��e�d�<�
�"�l�B݁�J��ƹF��Z�� ��b�%�u�h��0�(�������l��X�����e�
�
� �o�l����s���G��^\�� ��c�
�g�i�w�l�W����ο�T��������;� �
�g�4�(���&����U��[�����k�&�2�0��-��������9��G�����w�w�_�u�w�0�(������� R��N�U��u�=�;�}�>�3�Ǹ�&����gT��B��*���0�%��d�1��D���	�����Y�����:�&�
�#�o��^������D��N�����<�3�
�b��o�K���H�ƻ�V�D������-� ��9�(�(�������C9��1��*��
�g�u�u�>�3�ǿ�&����G9��V��0���0�&�u�e�l�}�WϪ�	����l��^�� ��c�
�g�i�w�l�W����Π�P9��]�� ��`�
�d�h�6�����&����lV�R��U��n�u�u�!�'�4����&����S��G\��H���w�"�0�u�;�>�!��&����R��GZ��U���6�;�!�9�o�m�W�������l�N�����<�<�
� �n�d����D������YN�����
�e�3�
�`��C������]��[��E���9�0�w�w�]�}�W���&����ZP��B1�@���u�h�w�w� �8�Wǲ�����9��hW�*��h�4�
�:�$�����I�Ʃ�@�L�U���!�%�<�<�>�n�(���A�ӓ�F�L�U���;�}�:�
��d����@ƹ��[��G1�����9�g�
�|�2�.�W��B�����h��*��� �b�l�%�w�`�U�������
��h8�� ��`�%�u�u�'�>�����ޓ�F��D��E��0�1�7�=�!�W