-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��a��c���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�4�0��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�^ �����
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W�������T��h��U���������!���6���F��@ ��U���_�u�u�;��3�������/��d:��9�������w�n�W������]ǻN�����;�0�b�0�c�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��a��R1�����o��u����>���<����N��
�����e�n�u�u�>�����&Ĺ��F��~ ��!�����
����_������\F��d��Uʼ�
�4�2�
���W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V �����!�:�
�g�2�m�Mϗ�Y����)��tUךU���;��;�4��3����H����F��~ ��!�����
����_������\F��d��Uʼ�
�4� �9�8�)����K����\��yN��1�����_�u�w�3�:�������G��h_����o��u����>���<����N��
�����e�n�u�u�>���������A	��\��*���u������4�ԜY�ƥ�l+��B�����:�
�g�0�b�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��~��V�����9�d�
�
�w�}�9ύ�=����z%��N�����4� �9�:�#�2�(������/��d:��9�������w�n�W������]ǻN�����<�&�a�0�g�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��t��D1����o��u����>���<����N��
�����e�n�u�u�>�����&ǹ��F��~ ��!�����
����_������\F��d��Uʼ�
�4�;�
���W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V��*ފ�
�u�u����;���:����g)��]����!�u�|�_�w�}��������l��T��;ʆ�������8���J�ƨ�D��^����u�;��<�$�i���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF��Y1�����a�0�b�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϷ�&����G9��N��U���
���n�w�}����/�ԓ�lV�'��&���������W��Y����G	�UךU���;��
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƥ�l6��1��G���u��
���(���-��� W��X����n�u�u�<���E���J����}F��s1��2������u�d�}�������9F���&���
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���*����V9��N��U���
���
��	�%���Hӂ��]��G�U���4�
�0� �9�m�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���R��R����o������0���/����aF�N�����u�|�_�u�w�-��������	F��cN��1��������}�D�������V�=N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӇ��A��E ��U��� �u��
���(���-��� W��X����n�u�u�4��8����L����f2��c*��:���
�����l��������l�N��*��� �;�c�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���	����F�� N�:���������4���Y����W	��C��\�ߊu�u�%�'�#�/�(���Y����`2��{!��6�����u�f�w�2����I��ƹF��G1�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}��������lW��N��!ʆ�������8���J�ƨ�D��^����u�%�'�!�%��F��6����g"��x)��*�����}�d�3�*����P���F��h��Oʜ�u��
���}�L����ƓR��^�����u�0�4�u�1�0�1��?�Ъ�9��N��U���u�6�;�!�9�}��������\��h_��U���
���u�j�z�P�ԜY�Ư�]��Y�����;�!�9�2�4�m�Mύ�=����z%�
N��R�ߊu�u�:�&�6�)����-����l ��h^��U���
���
��	�%���Kӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��Q��D��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��d�w�_�u�w�2����Ӈ��`2��C]�����u�u��
���(���-��� T��X����u�h�w�e�g�m�G��I����V��^�E��e�d�e�n�w�}��������R��c1��A���8�f�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�d�e�u�W�W�������]��G1��*���
�&�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�g�m�L���YӅ��@��CN��*���&�c�3�8�b�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�m�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�l�G��I��ƹF��X �����4�
��&�o�;���Cӵ��l*��~-��0����}�g�1� �)�W���C���V��^�E��e�e�e�e�g�m�F��I����l�N�����;�u�%���)�(���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��	���&����
F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����U��^��U���
���
��	�%���Kӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��h��*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��h��F���8�d�u�u���8���&����|4�\�����:�e�u�h�u�m�G��I����V��^�D��e�e�e�e�g�f�W�������R��V��!���d�
�&�
�d�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��d�e�e�e�g�m�G���s���P	��C��U����
�!�`�1�0�F���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�d�e�g�m�G��I���9F������!�4�
��$�l�(���&���5��h"��<������}�e�9� ���Y���F�^�E��e�e�e�e�f�m�G��I����V��d��Uʶ�;�!�;�u�'��(���N����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�F��I����V��^�W�ߊu�u�:�&�6�)����-����9��Z1�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��H����V��^�E��e�n�u�u�4�3����Y����g9��W�����m�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�w�]�}�W���
������d:�����3�8�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�g�
�&��m�Mύ�=����z%��r-��'���g�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%��
�!�e�;���Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
��.�E܁�
����\��c*��:���
�����o��������\�^�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-�$����ғ�@��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����GT��Q��G���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�*���
�`�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1��*���b�3�8�g�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�G��Y����\��V ������&�g�
�$��@��*����|!��h8��!���}�g�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%��
�#�d����K����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��	���&����_�=��*����
����u�EϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}����&����l ��h]�Oʆ�������8���J�ƨ�D��^��O���e�d�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������l��1����u�u��
���(���-��� T��X����u�h�w�d�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��c1��Fي�&�
�g�o���;���:����g)��]����!�u�|�o�w�l�G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�d�f�g�$���5����l0��c!��]���:�;�:�e�w�`�U���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�l�G��*����|!��h8��!���}�u�:�;�8�m�W��[����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������wF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EU��^��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�E���_�u�u�:�$�<�Ͽ�&����G9��\��D��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��d�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�d�w�_�w�}��������C9��Y����
�a�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�e�l�}�WϽ�����GF��h�����#�g�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�f�
�a�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�l�G��Y����\��V �����:�&�
�#�e�l�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��*��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�E���_�u�u�:�$�<�Ͽ�&����G9��\��3��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��d�n�u�u�4�3����Y����\��h��*���u��
����2���+����W	��C��\��u�e�e�n�w�}��������R��X ��*���g�g�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�D݁�8����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��H����]ǻN�����4�!�4�
�8�.�(���K�׉�	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>��������V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����R��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EP��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h]��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��Z��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��A]��A��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����\��h��A��o������!���6��� F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��d�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�e�w�]�}�W���
������T�����f�a�o����0���/����aF�
�����e�u�h�w�g��}���Y����G�������!�9�f�d�m��3���>����v%��eN��U���;�:�e�u�j��G���s���P	��C��U���6�;�!�9�e�o�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�d�1�"�#�}�^��Y����l�N�����;�u�%�6�9�)����?����`2��{!��6�����u�b�3�*����P���W��_�D��u�u�6�;�#�3�W�������l
��1�Oʆ�������8���K�ƨ�D��^��O���e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2����˹��	F��s1��2������u�`�9� ���Y���F�^�E��n�u�u�6�9�)����	����@��A_��A��u�u��
���(���-���R��X����u�h�w�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����\��c*��:���
�����i��������\�_�E��e�e�e�e�u�W�W�������]��G1�����9�d�
�e�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�N���u�6�;�!�9�}��������EW��^�Oʆ�������8���H�ƨ�D��^��O���e�e�e�d�g�m�G��B�����D��ʴ�
�:�&�
�!�h�C��Cӵ��l*��~-��0����}�a�1� �)�W���C���V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��Dڊ�u�u��
���(���-���
F��@ ��U���o�u�e�e�g�m�G���s���P	��C��U���6�;�!�9�f��1���Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���W��_�D��d�d�d�w�]�}�W���
������T�����d�
��o���;���:����g)��_����!�u�|�o�w�m�G��I����W��_�N���u�6�;�!�9�}��������EW��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(ؘ�I����\��c*��:���
�����l��������\�^�D��d�d�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������ES��T��!�����
����_�������V�S��E��d�n�u�u�4�3����Y����\��h��*���u��
����2���+����W	��C��\��u�e�e�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�l�G��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��I���9l�N�����u�%��
�$�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G��B�����E�����&�
�;�:�>�:�Mϭ�����9F������!�u�&�
�9�2�����ƭ�l%��Q��Oʦ�2�4�u�&�u�2���Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����W�,��9���n�u�u�&�0�<�W���L����l��h�����e�o�����4���:����W��X����n�u�u�&�0�<�W���L����l��h��U����
���l�}�Wϭ�����U��h]�*���
�e�o����0���/����aF�N�����u�|�_�u�w�4�������� V��R1�����0�&�u�u���8���&����|4�N�����u�|�_�u�w�4�������� V��R1����o������}���Y����R
��U1��F���0�e�"�d�m��3���>����F�D�����7�`�f�`�2�m����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*ߊ�e�
�
�
�3�/���Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*ߊ�e�
�
�
�2�}�W���&����p]ǻN�����9�3�
�
�g��(ށ�I����g"��x)��*�����}�d�3�*����P���F��P ��U���`�f�`�0�f�<����
����`2��{!��6�����u�d�3�*����P���F��P ��U���`�f�`�0�f�>�F��*����|!��d��Uʦ�2�4�u�7�b�n�B���H����\��c*��:���n�u�u�&�0�<�W���L����l��h
�Oʆ�������8���J�ƨ�D��^����u�<�;�9�1��(��&����R��R��U����
�����#���Q�ƨ�D��^����u�<�;�9�1��(��&����P��N��1�����_�u�w�4�������� V��R1�����u��
����2���+������Y��E��u�u�&�2�6�}����J�ӓ�lT��S
����o������!���6�����Y��E��u�u�&�2�6�}����J�ӓ�lT��R_��U���
���n�w�}�����ƪ�lS��[��*؊�0�u�u����>��Y����Z��[N��*ߊ�e�
�
�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��1�@ي�1�'�&�e�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƪ�lS��[����o������}���Y����R
��U1��D���
�e�o����0���/����aF�N�����u�|�_�u�w�4��������_��h�����d�o�����4���:����V��X����n�u�u�&�0�<�W���L���� 9��N�&������_�w�}����Ӏ��9��]�����u��
���f�W���
����_F��h[��L���1�u�u����>���<����N��
�����e�n�u�u�$�:��������V��h�����4�
� �g�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��B��*���
�1�'�2�'�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʷ�3�`�l�l�6�9�(���&����\��c*��:���
�����}�������9F������7�3�`�d�a���������F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�;�B��Oʹ��W��R	��A��o������!���6�����Y��E��u�u�&�2�6�}����H����R��h	��*���a�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӊ��9��V�����'�2�g�a�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������F ��h_�A���1�
�0�
�"�i�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�� ���
�m�a�4�3�����M���5��h"��<������}�w�2����I��ƹF��^	��ʼ�d�3�
�`�o�-�W���-����t/��a+��:���g�1�"�!�w�t�}���Y����R
��h_�����a�d�o����0���/����aF�
�����e�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��n�W���6����}]ǻN�����9�!�%�3��h�C���Y�Ɵ�w9��p'��#����u�c�u�8�3���B�����Y�����'�2�g�c�w�}�#���6����e#��x<��C���:�;�:�e�l�}�Wϭ�����V��T��@���
�`�g�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��X
�����
�d�
�
��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�;�1�
�2�0�E����ד�V��W�Oʆ�������8���Hӂ��]��G�U���&�2�4�u�'�.��������l��h��*���u��
���f�W���
����_F��h��*���
�`�u�u���6��Y����Z��[N�����;�a�3�
�b�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�l��h�����
�!�g�3�:�l�W���-����t/��=N��U���;�9�4�
�>�����O����q)��r/�����u�<�;�9�2�4����J����S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�'�.��������l��1����u�u��
���L���Yӕ��]��V�����1�
�l�u�w��;���B�����Y�����<�
�&�$���������� F��d:��9����_�u�u�>�3�Ͽ�&����Q��^�Oʗ����_�w�}����Ӈ��@��T��*���&�d�
�&��i�Mύ�=����z%��N�����4�u�%�&�0�?���@����|)��v �U���&�2�4�u��1�(���&����lW��Q��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϸ�&����\��X��DҊ�0�
�`�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�l��h�����
�!�b�3�:�l�W���-����t/��=N��U���;�9�4�
�>�����J����q)��r/�����u�<�;�9�#�-�E܁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��n����K����	F��s1��2������u�a�}�������9F������0�<�6�;�e�;�(��A����	F��s1��2������u�g�9� ���Y����F�D����� �
�
�`��m�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��G1�����0�
��&�f�����N����g"��x)��N���u�&�2�4�w�-��������R�,��9���n�u�u�&�0�<�W���&ƹ��_��N�&���������W��Y����G	�UךU���<�;�9�4��4�(�������@��h��*��o������}���Y����R
��G1�����1�f�c�o���2���s���@��V����� �d�e�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��O=�����
�b�'�2�e�i�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��U��@��f�
�
�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������D�����
��&�g��.�(��Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}����&����l��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�4���������C9��h��*���
�c�f�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�g�
�&��l�Mύ�=����z%��N�����4�u�%�&�0�?���A����|)��v �U���&�2�4�u�"��(��I����l��N��1��������}�D�������V�=N��U���;�9�6�
�#���������l��h��*��m�o�����4���:����U��S�����|�_�u�u�>�3�ϼ��ӓ�T��R1�����u��
����2���+������Y��E��u�u�&�2�6�}����&����	��h\�����'�2�g�e�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��r"��!���
�c�3�
�a�k����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����� �
�a�/���H����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʡ�%�a�
� �f�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
�0�
�b�o�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��V�� ��f�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����^��R	��B��o������!���6�����Y��E��u�u�&�2�6�}��������Z9��h_�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��R	��B��o������!���6�����Y��E��u�u�&�2�6�}��������Z9��h_�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��R	��B���o������!���6�����Y��E��u�u�&�2�6�}��������Z9��h_�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��R	��B��o������!���6�����Y��E��u�u�&�2�6�}��������Z9��h_�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��R	��B��o������!���6�����Y��E��u�u�&�2�6�}�$���=����G9��h��*��f�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�&����P��h=����
�&�
�g�m��3���>����F�D�����%�&�2�7�3�i�N��;����r(��N�����4�u�'�
�"�l�Fہ�K����g"��x)��*�����}�d�3�*����P���F��P ��U���6�
�m�'�0�o�B���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����g��!�o��(���K����CU�=��*����
����u�FϺ�����O��N�����4�u��-��	����&�ғ�l��h\�A��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���&����\��c*��:���
�����}�������9F������6�
� ���8���&����U��Z�����u��
����2���+������Y��E��u�u�&�2�6�}����7����V��V��*؊�0�
�b�a�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�g�
�$��D��*����|!��d��Uʦ�2�4�u�%�$�:����M���$��{+��N���u�&�2�4�w�����-����l+��C����
�0�
�b�b�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h[��F���0�e�$�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ư�l
��q��9���
�f�0�e�%�:�E��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����<�
�&�$����������F��d:��9����_�u�u�>�3�Ͽ�&����Q��Y�Oʗ����_�w�}����Ӗ��G��^1��*��m�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����^��h��*��e�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�&����P��h=����
�&�
�`�m��3���>����F�D�����%�&�2�7�3�i�O��;����r(��N�����4�u�!�`�f�e�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&������!�%��B�������F��d:��9�������w�n�W������]ǻN�����9�4�
�<��.����&����l ��h\�Oʆ�����]�}�W�������C9��P1����l�o�����}���Y����R
��C1��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������w#��e<�����b�'�2�g�f�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h[��M���0�e�$�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ư�l/��r6��'���8�d�e�0�g�/���K����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʹ�
�
�m�c�2�l����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*������0�:�l�G���H����lT��N�&���������W��Y����G	�UךU���<�;�9�9���O����֓�F��d:��9�������w�n�W������]ǻN�����9�6�
����%�������l��h��*��c�o�����4���:����U��S�����|�_�u�u�>�3�ϲ�&ƹ��P��h_��D��������4���Y����W	��C��\�ߊu�u�<�;�;�>�(���<����G��h_�*���
�0�
�m�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��~ ��-���!�'�
�l�%�:�E��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����<�
�&�$����������F��d:��9����_�u�u�>�3�Ͽ�&����Q��]�Oʗ����_�w�}����Ӏ��z(��o/�����
�d�'�2�e�j�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��T��;�����0�8�f�i��������Q��N��1��������}�D�������V�=N��U���;�9�6�
���6�������R��h_�����m�d�o����0���/����aF�N�����u�|�_�u�w�4��������w#��e<�����`�
�
�
�2��O��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��������!�%��Bف�&¹��T9��_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�����@ǹ��\��c*��:���
�����}�������9F������<�f�'�2�e�d�W���-����t/��a+��:���g�1�"�!�w�t�}���Y����R
��G1�����0�
��&�d�����@����g"��x)��N���u�&�2�4�w�-��������S�,��9���n�u�u�&�0�<�W���&�֓�F9��^��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����_��T��!�����
����_������\F��d��Uʦ�2�4�u�-�#�2�ށ�����9��T��!�����
����_�������V�=N��U���;�9�<�a�1��E���	����`2��{!��6�����u�d�3�*����P���F��P ��U���
�0�
�l�n�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��^	������
�!�g�1�0�D���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�)���&����W��G_��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�:��F�������F��d:��9�������w�k�W������]ǻN�����9�0�<�6�9����IĹ��\��c*��:���
�����}�������9F������7�3�`�f�b�8�G�������F��d:��9�������w�l��������l�N�����u� �
�
�g��(߁�����`2��{!��6�ߊu�u�<�;�;�?����J�ӓ�lV��N�&���������W��Y����G	�UךU���<�;�9�7�1�h�D����֓�W��D�Oʆ�������8���Hӂ��]��G�U���&�2�4�u�"��(��&����P��N��1�����_�u�w�4��������lU��h��*���u�u��
���L���Yӕ��]��U��@��`�0�e�1�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Q��1�@���d�4�1�0�$�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[��Eߊ�
�
�0�u�w�	�(���0��ƹF��^	��ʷ�3�`�f�`�2�l����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����f�`�0�d�6�9����Y�Ɵ�w9��p'��#����u�d�1� �)�W���s���@��V�� ���
�e�
�
��8�W���-����t/��=N��U���;�9�7�3�b�n�B���H����\��c*��:���n�u�u�&�0�<�W���&ƹ��9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�(�(ځ�Iƹ��9��S�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�?����J�ӓ�lT��R^��U���
���n�w�}�����Ʈ�U9��^�����$�u�u����>���<����N��
�����e�n�u�u�$�:�������� V��R1�����0�&�u�u���8���&����|4�N�����u�|�_�u�w�4��������lU��h��*���u�u��
���L���Yӕ��]��U��@��`�0�g�"�f�g�$���5����l�N�����u� �
�
�g��(݁�H����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�`�
�3�/���Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����l�l�6�e�m��3���>����F�D����� �
�
�`��9����H����g"��x)��*�����}�u�8�3���B�����Y�����`�l�l�6�f�g�$���5����l�N�����u� �
�
�b�����Y����)��tUךU���<�;�9�7�1�h�N�������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʷ�3�`�d�c��9����I����g"��x)��*�����}�u�8�3���B�����Y�����`�d�c�
�2�}�W���&����p]ǻN�����9�7�3�`�f�k�(�������\��c*��:���
�����}�������9F������7�3�`�d�a�����Y����)��tUךU���<�;�9�7�1�h�F��&����	F��s1��2���_�u�u�<�9�1����L����
9��T��!�����
����_������\F��d��Uʦ�2�4�u� ���N����֓�W��D�Oʆ�������8���Hӂ��]��G�U���&�2�4�u�"��(��H����l��T��!�����n�u�w�.����Y����9��_��*ڊ�e�o�����4���:����V��X����n�u�u�&�0�<�W���&ƹ�� W��h^�����&�d�o����0���/����aF�
�����e�n�u�u�$�:��������_��h��*���u�u��
���L���Yӕ��]��U��@��f�
�
�
�2�}�W���&����p]ǻN�����9�7�3�`�e�n�(���&���5��h"��<������}�w�2����I��ƹF��^	��ʷ�3�`�g�f���(�������\��c*��:���
�����}�������9F������7�3�`�g�d��(ށ�����`2��{!��6�ߊu�u�<�;�;�?����K����V9��F^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�"��(��H����l��E��D��������4���Y����\��XN�N���u�&�2�4�w�(�(ځ�@�ד�lW��R_��U���
���n�w�}�����Ʈ�U9��W�*���
�0�u�u���8���B�����Y�����`�g�f�
���F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*ߊ�c�e�0�e�6�9����Y�Ɵ�w9��p'��#����u�d�1� �)�W���s���@��V�� ���
�c�e�0�g�>�G��*����|!��d��Uʦ�2�4�u� ���A����֓�W��D�Oʆ�������8���Hӂ��]��G�U���&�2�4�u�"��(��I����l��T��!�����n�u�w�.����Y����9��^��*ڊ�0�u�u����>��Y����Z��[N�����d�g�
�
��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��B��*��e�0�d�4�3�8����Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T����*ߊ�c�e�0�d�4�m�Mύ�=����z%��N�����4�u� �
��k�G���H����A��N�&���������W������\F��d��Uʦ�2�4�u� ���A����ד�VW�=��*����n�u�u�$�:��������P��h��*���u�u��
���L���Yӕ��]��U��@��g�
�
�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h[��Dڊ�
�
�1�'�$�m�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Q1��L���0�e�6�e�m��3���>����F�D����� �
�
�d���(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�� ���
�d�
�
��9����H����g"��x)��*�����}�u�8�3���B�����Y�����`�l�e�0�g�>�F��*����|!��d��Uʦ�2�4�u� ���F߁�&ù��F��d:��9����_�u�u�>�3�ϼ��ӓ�V��h^��D��������4���Y����W	��C��\�ߊu�u�<�;�;�?����@�֓�lW��S
����o������!���6�����Y��E��u�u�&�2�6�}����&����V9��T�Oʆ�����]�}�W�������F ��hW�*���
�e�o����0���/����aF�N�����u�|�_�u�w�4��������l_��h��*���'�&�d�o���;���:����g)��_�����:�e�n�u�w�.����Y����9��1��D���d�o�����4�ԜY�ƿ�T����*ߊ�d�
�
�
�2�}�W���&����p]ǻN�����9�7�3�`�n�m��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʷ�3�`�d�f���(�������\��c*��:���
�����}�������9F������7�3�`�d�d��(߁�����`2��{!��6�ߊu�u�<�;�;�?����H����V9��V
�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����L���� 9��1��D�������W�W���������h[��F���0�e�"�d�m��3���>����F�D����� �
�
�f�d�8�G���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����`�d�f�
������
���5��h"��<������}�w�2����I��ƹF��^	��ʷ�3�`�d�f���(���Y�Ɵ�w9��p'�����u�<�;�9�5�;�B��J����9��S�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�?����H����V9��T�Oʆ�����]�}�W�������F ��h_�F���d�"�d�o���;���:���F��P ��U���
�
�f�f�2�l����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����d�f�
�
��9����I����g"��x)��*�����}�u�8�3���B�����Y�����`�d�f�
������Y����)��tUךU���<�;�9�7�1�h�F��&����R��R��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�;�B��J����9��N�&������_�w�}����ӄ��lS��]�����"�d�o����0���s���@��V�� ���
�f�f�0�e�9�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��[��*��m�4�1�0�$�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������
��1�MҊ�0�u�u����>��Y����Z��[N��*ߊ�c�m�4�1�2�.�W���-����t/��a+��:���d�1�"�!�w�t�}���Y����R
��C1��D��
�0�u�u���8���B�����Y�����
�c�m�"�f�g�$���5����l�N�����u�!�`�d�o��F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����@��a�
�
�
�3�/���Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*ߊ�m�c�0�e�4�m�Mύ�=����z%��N�����4�u�!�`�f�i�(���&����V��T��!�����
����_�������V�=N��U���;�9�9�
��e�A���I����\��c*��:���n�u�u�&�0�<�W���L����9��1��D�������W�W�������
��1�A܊�
�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӊ��9��X��*ۊ�1�'�&�e�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ơ�lS��Z�����6�e�o����0���s���@��V�����d�a�
�
��9����H����g"��x)��*�����}�u�8�3���B�����Y�����
�m�c�0�f�>�F��*����|!��d��Uʦ�2�4�u�!�b�l�Cف�&¹��F��d:��9����_�u�u�>�3�ϲ�&ƹ��P��h_��D��������4���Y����W	��C��\�ߊu�u�<�;�;�1�(ځ�O�ӓ�lV��S
����o������!���6�����Y��E��u�u�&�2�6�}����L����V9��T�Oʆ�����]�}�W�������G9��X�*���
�e�o����0���/����aF�N�����u�|�_�u�w�4��������P��h��*���'�&�d�o���;���:����g)��_�����:�e�n�u�w�.����Y����lS��1��E���d�o�����4�ԜY�ƿ�T����@���l�
�
�
�2�}�W���&����p]ǻN�����9�9�
�
�a�h��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʹ�
�
�c�`�2�l��������	F��s1��2������u�f�9� ���Y����F�D�����!�`�`�l���(���Y�Ɵ�w9��p'�����u�<�;�9�;��(��L����l��N��1��������}�D�������V�=N��U���;�9�9�
��k�B���H����A��N�&���������W������\F��d��Uʦ�2�4�u�!�b�h�Nځ�&¹��F��d:��9����_�u�u�>�3�ϲ�&ƹ��
S��h_�����u��
���f�W���
����_F��h[��C���0�d�1�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ơ�lS��W�����4�1�0�&�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������G9��X�*���
�0�u�u���8���B�����Y�����
�c�`�0�e�,�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��[��*��`�0�g�4�3�8����Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T����@���l�
�
�
�2�}�W���&����p]ǻN�����9�9�
�
�a�h�������5��h"��<��u�u�&�2�6�}����L����V9��S_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�"��(��M����A��N�&���������W������\F��d��Uʦ�2�4�u� ���O������5��h"��<��u�u�&�2�6�}����&����l��N��1��������}�D�������V�=N��U���;�9�7�3�b�l�Oہ�����@W�=��*����
����u�W������]ǻN�����9�7�3�`�f�e�(���Y�Ɵ�w9��p'�����u�<�;�9�5�;�B��Aǹ��F��d:��9����_�u�u�>�3�ϼ��ӓ�^��S_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��8�(��A����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$���܁�
����	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������\��C��*��
�
�0�
�c�d�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��*���$��
�!��.�(���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����l5��D�����b�o�����4�ԜY�ƿ�T�������7�1�m�m�m��8���7���F��P ��U���'�2�d�c�w�}�#���6����e#��x<��Gʱ�"�!�u�|�]�}�W�������C9��P1������&�d�
�$��G��*����|!��d��Uʦ�2�4�u�%�$�:����A���$��{+��N���u�&�2�4�w���������\��h��*��g�o�����4���:����T��X����n�u�u�&�0�<�W���
����@��d:�����3�8�d�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��h�W���6����}]ǻN�����9�4�
�<��.����&����l ��h\�Oʆ�����]�}�W�������C9��P1����l�o�����}���Y����R
��1����m�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�&����P��h=����
�&�
�e�m��3���>����F�D�����%�&�2�7�3�e�N��;����r(��N�����4�u�f�'�0�l�N���Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T�������6�0�
��$�n�(���&���5��h"��<��u�u�&�2�6�}��������l^��T��:����n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��d�W���6����}]ǻN�����9�4�
�<��.����&����U��N�&������_�w�}����Ӈ��@��U
��L��o�����W�W���������h�� ��b�
�d�o���;���:����g)��X����!�u�|�_�w�}����Ӓ��lT��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�4�
�<��.����&����l ��hW��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��G1�*���d�e�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������A��B1�Eߊ�e�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����S��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-����L�ғ�F��d:��9�������w�n�W������]ǻN�����9�2�%�3��h�C���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�
�`�l�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��*���l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����V��B1�BҊ�g�o�����4���:����W��X����n�u�u�&�0�<�W����ԓ�l ��X�*��o������!���6���F��@ ��U���_�u�u�<�9�1����/�ԓ�F9��_��A��������4���Y����\��XN�N���u�&�2�4�w�2�(���&����S��G_��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�:��(�������P��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��(���&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�&����Q��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�8��(ہ�����9��T��!�����
����_�������V�=N��U���;�9�9�6��h����O�ѓ�F��d:��9�������w�o�W������]ǻN�����9�!�%�<�>��(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�d�>�4�(�������9��T��!�����
����_�������V�=N��U���;�9�%��;��(���H����CW�=��*����
����u�FϺ�����O��N�����4�u�:�
�����H����\��c*��:���
�����}�������9F������9�6��b�1��@���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʡ�%�<�<�
��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�d�<�<�����J����\��c*��:���
�����}�������9F������;�!�=�d�1��@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���9�&�
� �f�i�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����g�3�
�b�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��X��؊� �d�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��V�� ��`�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����_��B1�Bߊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�֓�F9��_��G��������4���Y����\��XN�N���u�&�2�4�w�/�(���H����CT�=��*����
����u�W������]ǻN�����9�;�!�=�d�;�(��@����	F��s1��2������u�g�9� ���Y����F�D�����:�9�&�
�"�l�N܁�K����g"��x)��*�����}�u�8�3���B�����Y�����f�
� �d�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Fߊ� �d�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��X�� ��g�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����U��B1�Fڊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�ѓ�F9��[��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������T��^1��*��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��Z�����
� �d�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G_�� ��a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y���� P��R�����<�3�
�c�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��F���
�b�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���0�:�2�;�1��O���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�b�3�
�o�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
�
� �f�h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�l�<�3��e�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�
�
�8����NĹ��\��c*��:���
�����}�������9F������!�%�a�
�"�l�Eց�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�m�<�1��O���	����`2��{!��6�����u�e�3�*����P���F��P ��U��� ����#�/�(�������W��N�&���������W��Y����G	�UךU���<�;�9�9�4�����@�ӓ�F��d:��9�������w�j��������l�N�����u�:�
�
��(�F��&���5��h"��<������}�e�9� ���Y����F�D�����8�
�
�
�����Kƹ��\��c*��:���
�����}�������9F������!�%�<�<�>�;�(��@����	F��s1��2������u�g�9� ���Y����F�D�����0�
�
�
��(�F��&���5��h"��<������}�c�9� ���Y����F�D�����8�
�
�
�����Jʹ��\��c*��:���
�����}�������9F������&�9�!�%�����O¹��\��c*��:���
�����}�������9F������&�9�!�%�����OĹ��\��c*��:���
�����}�������9F������'�!�g�<�>�4����&����l ��W�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l ��W�*��o������!���6���F��@ ��U���_�u�u�<�9�1����
����@9��h_�D���u�u��
���(���-���Q��X����n�u�u�&�0�<�W���������C1�*���0�%��d�1��N���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʡ�%�<�3�
�n�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���<�3�
�e�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��L���
�e�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��h��G��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����M����V��h�Oʆ�������8���Nӂ��]��G�U���&�2�4�u��l�F�������V��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-�Eׁ�&����R��G]��U���
���
��	�%���Iӂ��]��G�U���&�2�4�u��8����H¹��lT��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����-����G9��h�����%�
� �d�`��D��*����|!��h8��!���}�a�1�"�#�}�^�ԜY�ƿ�T����*���c�<�3�
�g�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���b�<�3�
�g�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���m�<�3�
�g�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��������;� �
�c�;�(��H����	F��s1��2������u�d�}�������9F������;�!�=�
�"�o�Nށ�K����g"��x)��*�����}�u�8�3���B�����Y�����g�
� �g�n��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��A܊� �g�e�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����U5��R��*��
�
� �g�e��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������d�d�g�d�1��F���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʦ�9�!�%�d�>�;�(��L����	F��s1��2������u�d�}�������9F������&�9�!�%�g�4����H�ԓ� F��d:��9�������w�n�W������]ǻN�����9�&�9�!�'�d����&����l��N��1��������}�D�������V�=N��U���;�9�3�
���#���&����U��[�����u��
����2���+������Y��E��u�u�&�2�6�}��������Z9��h\�A���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����9��Q��D���%�u�u����>���<����N��
�����e�n�u�u�$�:��������CU��^1��*��`�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U��^�����1�u�u����>���<����N��S�����|�_�u�u�>�3�Ϲ�	����S��h��Oʆ�����]�}�W�������C9��P1������&�d�
�$��O��*����|!��d��Uʦ�2�4�u�%�$�:����H����	F��x"��;�ߊu�u�<�;�;�:����&����l	��X
��Oʆ�������8���Mӂ��]��G�U���&�2�4�u�:��A���&����l	��X
��Oʆ�������8���Mӂ��]��G�U���&�2�4�u�:��D���&����l	��X
��Oʆ�������8���Mӂ��]��G�U���&�2�4�u�:��@���&����l	��X
��Oʆ�������8���Mӂ��]��G�U���&�2�4�u�'��(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����<�
�1�
�n�h�MϜ�6����l�N�����u�%�&�2�5�9�F��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����\��x!��4��u�u�&�2�6�}��������lW��T��:����n�_�u�w�2�����ơ�uP��q_��*ڊ�4�1�&�7�d�3�(���
���� 9��[������u�u�2�9�/����Y���F��sN�<�����_�u�w�}�W���&����vF��~ ��2���_�u�u�u�w�4�G���=���/��r)��N���u�u�u�1�9��>���Y�ƅ�g#��eUךU���u�u�:�!� ��?��0����v4�d��Uʥ�'�u�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�%�.���0�Ɵ�w9��p'�����u�u�u�<�g�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Y�����N�<����
�����#���Q����\��XN�N���u�u�u�:�4�9�W���7ӵ��l*��~-��0����}�u�:�9�2�G��Y���F��RN�<����
���l�}�W���Yӂ��GF��x;��&���������W��Y����G	�N����u�;�u�:�'�3���s�����G������c�e�d�1�m����&�Ԣ�lU��D1�*ۊ�4�
�&�u��}�WϹ�����NǻN��U����o�����}���Y���}3��d:��0������]�}�W���Y����l1��c&��U�����n�u�w�}�WϺ�¹��w2��N��!����_�u�u�w�}����.����\��y:��0���n�u�u�%�%�}�}���Y���W��T��;ʆ�������8���J�ƨ�D��^����u�u�u�<�f�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Y�����CN�:���������4���Y����W	��C��\���_�u�u�;�w�2������Ɠ9F������;�u��c�g�l�������� T��h]�����d��_�u�w�8����Y���F�N��U������n�w�}�W���7����g'��T��;����n�u�u�w�}����&����{F��~ ��2���_�u�u�u�w�4�F���=���/��r)��N���u�u�u�1�"��>���Y�ƅ�g#��eN����u�:�!�}�w�}�W�������	F��=��*����
����u�FϺ�����O��N��U���1�;�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����W�'��&���������W������\F��d��U���u�1� �u�w��W���&����p9��t:��U��1�"�!�u�~�t�}���Y����P	��X ���ߠ_�u�u�:�'�3����8����uW��h^��*ߊ�7�`�f�`�2�m�>�ԜY�ƫ�]��TN��U���u�u��!� �9���0����v4��N��U����1�0�&�6�:�W���7����a]ǻN��U���1�'�&��3�5�Mϗ�-����O��N�����u�_�u�u�w�}����Y����g"��x)��N���u�u�u�'�$�)�Mϗ�Y����)��tUךU���u�u�1�'�$�m�Mϗ�Y����)��t1��6���u�d�1�"�#�}�^�ԜY���F��N�<����
���l�}�W���Yӗ��	F��cN��1��������}�D�������V�=N��U���u�1�'�&�f�g�>���-����t/��a+��:���d�1�"�!�w�t�}���Y���P��N��U���
���n�w�}�W������/��d:��9����_�u�u�w�}�F��0�Ɵ�w9��p'��#����u�f�u�8�3���Y��ƹF��Y
�����;�;�n�_�w�}����������Z��Dܳ�e�3�`�3���N��0���F��Y�����u�u�u�u��)� �������}2��r<�U���u�u��1�2�.����Y�ƅ�g#��eUךU���u�u�1�'�$�
����Cӯ��v!��G�U���%�'�u�_�w�}�W�������z(��c*��:���n�u�u�u�w�/����Cӯ��`2��{!��6�ߊu�u�u�u�3�/���Cӯ��`2��{!��6�����u�e�3�*����P���F�N��E���u��
���L���Y�����N��!ʆ�������8���J�ƨ�D��^����u�u�u�1�%�.�F��0�Ɵ�w9��p'��#����u�e�1� �)�W���s���F�T�Oʜ�u��
���f�W���Y����VW�'��&������_�w�}�W���H����}F��s1��2������u�d�}�������]ǻN�����:�%�;�;�l�W�W�������]����C���d�3�e�3�b�?����J�ӓ�lV��dd��Uʲ�;�'�6�}�w�}�W���=����Z��T��;����n�u�u�w�}�6�������]��N��!����_�u�u�w�}����
����G�'��0���u�n�u�u�'�/�W�ԜY���F��\N�<����
���l�}�W���YӔ��V�'��&������_�w�}�W�������@V�'��&���������W������\F��d��U���u�6�e�o��}�#���6����9F�N��U��o������0���/����aF�N�����u�|�_�u�w�}�W�������\��yN��1��������}�FϺ�����O��N��U���6�d�o��w�	�(���0��ƹF�N�����u������4�ԜY���F��T��;ʆ�������8���J�ƨ�D��^��\�ߊu�u�;�u�8�-����B��ƹF��X�����u��c�e�f�;�G���L����lS��]�����_�u�u�2�8����s���F�s��"���=�o�����}���Y���r��R�����u�u����f�W���Y����W��D�����o�����t�}���Y����NǻN��U���9�u�u����;���:���F�N�����o��u����>��Y���F��S
����o��u����>���<����N��S�����|�_�u�u�w�}����Y����g"��x)��N���u�u�u�$�w�}�"���-����t/��a+��:���e�1�"�!�w�t�}���Y���R��R��U���������!���6�����Y��E��u�u�u�u�4�l�Mϗ�Y����)��tUךU���u�u�0�u�w��$���5����l�N��Uʱ�u�u�����0���/����aF�
�����e�u�n�u�w�8�Ͻ�����]��=d��Uʶ�8�:�0�!�:��Cߘ�O����U9��[��*��m��_�u�w�8����Y���F�N�����1�=�o����%�ԜY���F��S�����2�u�u����L���Y���'��E��"���=�o�����^�ԜY�Ƽ�A�=N��U���u�9�u�u���3���>����F�N�����!�o��u���8���B���F������e�o��u���8���&����|4�N�����u�|�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�&�}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y���F��S
����o��u����>���<����N��S�����|�_�u�u�w�}����Y����g"��x)��N���u�u�u�"�f�g�>���-����t/��=N��U���u�d�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������|3��d:��9�������w�n�W������F�=N��U���u�:�%�;�9�f�}���YӅ��C	��Y��4��e�d�3�e�1�h����L����F��=N��U���0�<�u�_�w�}�W�������W��N��!����_�u�u�w�}����
����T�'��0���n�u�u�u�w�����
����[F��~ ��2���|�_�u�u�8�)�_���Y�����T��;ʆ�����]�}�W���Y����GF��~ ��!�����n�u�w�}�WϿ�����F��~ ��!�����
����_�������V�=N��U���u�0�u�u���3���>����F�N�����u� �u����>���<����N��
�����e�n�u�u�w�}��������	F��=��*����
����u�W������]ǻN��U���0�u�u����;���:���F�N��D���u��
���L���Y�����N��U���
���
��	�%���Hӂ��]��G��N���u�0�1�6�:�2����s����V��=N��U���`�f�`�0�g��MϽ�����]��v(�E��3�e�3�`�1��(��&����F�P�����8�%�}�u�w�}�WϚ�����G�	N�Y���u�u�u��3�8�������R�N��U����1�0�&�>�)�W���K���F��E�����_�u�u�u�w�1�W�������XJǻN��U���0�0�u�k�6����Y���F��S
����h�u�7�`�d�h��������@��=N��U���u�0�u�k�1��(��&����P��=N��U���u�e�h�u�5�h�D����֓�JǻN��U���1�'�&�d�j�}����J�ӓ�lV��S
����_�u�u�u�w�8�W������� V��R1����_�u�u�u�w�8�W������� V��R1����_�u�u�u�w�l�J����ӓ�S��h^��D��_�u�u�7�b�n�B���H�����G������c�e�d�1�m�������� V��R1�U���2�;�'�6�:�-�_���Y���"��V9�����k�f�y�u�w�}�Wϟ�����a��RN��U���u�u�u�u��9��������X�d��Uʥ�'�u�4�u�]�}�W���Y����X��G1���ߊu�u�u�u�2�8�W�������GJǻN��U���1�'�&�e�j�}����J�ӓ�lW��S
����_�u�u�u�w�8�W������� V��R1����_�u�u�u�w�m�J����ӓ�S��h_��E�ߊu�u�u�u�3�/���D�ƪ�lS��[��*ۊ�1�'�&�d�]�}�W���Y����X��U1��F���0�d�6�d�]�}�W���Y����X��U1��F���0�d�"�d�]�}�W���Y���F��h[��Eߊ�
�
�d�n�]�}�W���L����l��h;��U���%�;�;�u��k�G���֓�lS��U1��F���0�e�u�u�0�3�������9F�N��U���4�<�!�u�i�n�[���Y���'��E��'���0�h�u�y�w�}�W���8����@��S��H���|�u�u�%�%�}����s���F�T��H���%�6�>�_�w�}�W�������X��G1���ߊu�u�u�u�3�/���D�ƪ�lS��[��*؊�1�'�&�e�]�}�W���Y����X��U1��F���0�g�6�e�]�}�W���Y���F��h[��Eߊ�
�
�e�_�w�}�W�������@W�	N��*ߊ�e�
�
�
�3�/���s���F�T�H���7�`�f�`�2�o���s���F�@�H���7�`�f�`�2�o� ��s���F�S_��Kʳ�
�
�e�
���F��s���U��h_�F���o�6�8�:�2�)����Mà��U9��Q1�����
�l�f�u�w�:����Ӌ��NǻN��U���4�4�<�!�w�c�D��Y���F��S
�����;�0�h�u�{�}�W���Yӧ��A��`����u�|�u�u�'�/�W���Y���F�N����u�%�6�>�]�}�W���Y����GF������_�u�u�u�w�9����I���U��h_�F���1�0�&�y�w�}�W������F��h[��L���6�e�_�u�w�}�W��D�ƪ�lS��[�����u�u�u�u�6�9����Y����Q9��W�*���'�&�d�_�w�}�W������ ��1�@ي�0�y�u�u�w�}� ��D�ƪ�lS��[����_�u�u�u�w�l�J����ӓ�
S��S_����u�7�3�`�d�h����,����\��Y��U���c�e�d�3�g�;�B����ӓ�S��h^ךU���0�0�<�u�6�}�}���Y���w��`����u�g�_�u�w�}�W�������R��S�A�ߊu�u�u�u�3�/�������F��=N��U���!�8�%�}�w�}�W������F��h��Y���u�u�u�'�$�)�J���	����l�N��Uʴ�1�0�&�u�i�?����J�ӓ�lV��S
����_�u�u�u�w�8�W�������lU��h��*���y�u�u�u�w�,�W�������lU��h��*��_�u�u�u�w�9����H���Q��1�@���e�4�1�0�$�q�W���Y����VW�	N�����f�`�0�e�4�l�}���Y���D��
P�� ���
�e�
�
��8�[���Y�����
P�� ���
�e�
�
��l�L�ԜY�Ʈ�U9��^����� �o�6�8�8�8�ϳ�?����P��1��@���3�`�f�`�2�m�W�������Z��V�����u�u�u�4�6�4����G����9F�N��U���'�&��;�2�`�W��Y���F��S
�����1�=�h�u�~�}�WϮ��ơ�CF�N��U���6�>�h�u�'�>��ԜY���F��D��H���%�'�!�_�w�}�W�������@V�	N�����f�`�0�d�6�9����U���F���U��7�3�`�f�b�8�F���I���F�N��U��7�3�`�f�b�8�F���U���F������d�h�u� ���Gځ�&¹��W��D_�U���u�u�6�d�j�}����&����V9��T����u�u�u�0�w�c����L����l��h��Y���u�u�u�1�w�c����L����l��h
�N�ߊu�u� �
��m�(���&����P	��X ��ʸ��a��c���(ځ����� V��R1�U���2�;�'�6�:�-�_���Y���"��V9�����k�f�y�u�w�}�Wϟ�����a��RN��U���u�u�u�u��9��������X�d��Uʥ�'�u�4�u�]�}�W���Y����X��G1���ߊu�u�u�u�2�8�W�������GJǻN��U���1�'�&�e�j�}����&����V9��V
�����y�u�u�u�w�>�G��Y����9��1��G���e�_�u�u�w�}�G��Y����9��1��G���y�u�u�u�w�<����
�����h[��Eߊ�
�
�1�'�$�l�}���Y���P��
P�� ���
�e�
�
��8�[���Y�����S����`�f�`�0�e�*�F�ԜY���F��S����`�f�`�0�e�9�^�ԶY����F ��hW�*���u�:�%�;�9�}�6��I����lV��h[�� ���
�e�
�
�]�}�W�������^��d��U���u��!��3�5�J���K���F�N�����&�4�2�u�i�i�}���Y���r��R�����u�k�g�_�w�}�������9F�N��U���u�k�4�
�;�q�W���Y����V��S����&�y�u�u�w�}��������X��B��*���
�1�'�&�g�W�W���Y�Ư�F���*ߊ�`�
�0�y�w�}�W��������h[��@ӊ�e�_�u�u�w�}����
���F��Q1��L���4�1�0�&�{�}�W���YӅ��[�U��@��l�6�d�_�w�}�W��������h[��@ӊ�0�y�u�u�w�}����Gӄ��lS��W��D��_�u�u� ���B���,����\��Y��U���c�e�d�3�g�;�B����ӓ�S��h^ךU���0�0�<�u�6�}�}���Y���w��`����u�g�_�u�w�}�W�������R��S�A�ߊu�u�u�u�3�/�������F��=N��U���!�8�%�}�w�}�W������F��h��Y���u�u�u�'�$�)�J���	����l�N��Uʴ�1�0�&�u�i�?����H����R��R��Y���u�u�u�6�g�`�W���&ƹ��_��R^�U���u�u�$�u�i�?����H����BV�N��U���4�1�0�&�w�c����L����
9��S�����u�u�u�u�4�l�J�������S��h��Y���u�u�u�"�f�`�W���&ƹ��_��R_�U���u�u�1�u�i�?����H����WW�=d��Uʷ�3�`�g�f���(���Y����\��CN��3���c�
�
������&����l��=N��U���0�<�u�4�w�W�W���Y�ƈ�G��S��H���y�u�u�u�w�����
����VF�Z�U���u�u��1�2�.����Y���l�N�����4�u�_�u�w�}�W���Y����C9��\BךU���u�u�0�0�w�c����
��ƹF�N�����&�e�h�u�"��(��H����l��E��E�ߊu�u�u�u�2�}�Iϼ��ӓ�
U��R1����_�u�u�u�w�m�J�������_��h��*��_�u�u�u�w�9����H���Q��1�Fۊ�
�
�1�'�$�l�}���Y���P��
P�� ���
�l�d�0�g�>�F�ԜY���F��N��U���
�
�l�d�2�m� ��s���F�S_��Kʷ�3�`�g�f���(��B���F��Q1��G��
�
�
�u�w�2�����ơ�uP��q_��*ڊ�
�
� �
��m�(���s���T��E�����}�u�u�u�w��������F��d��U���u��1�0�$�<����G����F�N��4���0�&�<�!�w�c�E�ԜY�Ƽ�A��V�����u�u�u�9�w�c������ƹF�N�����u�k�4�
�$�q�W���Y����W��D�H��� �
�
�l�f�8�F�������JǻN��U���0�u�k�7�1�h�E��&����P��=N��U���u�e�h�u�"��(��H����l��=N��U���u�1�'�&�f�`�W���&ƹ�� W��h_�����&�d�_�u�w�}�W���Y����F ��h\�D���d�6�d�_�w�}�W��������h[��L���0�d�"�d�]�}�W���Y���F��Q1��G��
�
�
�d�l�W�W�������P��h��*���u�:�%�;�9�}�6��I����lV��h[�� ���
�e�
�
�]�}�W�������^��d��U���u��!��3�5�J���K���F�N�����&�4�2�u�i�i�}���Y���r��R�����u�k�g�_�w�}�������9F�N��U���u�k�4�
�;�q�W���Y����V��S����&�y�u�u�w�}��������X��B��*��e�0�e�4�3�8���Y���F��R^��Kʷ�3�`�d�g���(���U���F��H��� �
�
�c�g�8�G���U���F������d�h�u� ���A����֓�W��D����u�u�u�0�w�c����L����9��1��D�ߊu�u�u�u�2�}�Iϼ��ӓ�T��R1����_�u�u�u�w�l�J�������P��h��*��n�_�u�u�"��(��I����l3������;�u��c�g�l�����ӓ�F ��h]�*���_�u�u�0�2�4�W���Y���F�N�����1�=�h�u�e�W�W���Y�ƍ�W��D<�����k�a�_�u�w�}�W�������Z��S�G�ߊu�u�:�!�:�-�_���Y�����S����9�y�u�u�w�}�������R��D�U���u�u�4�1�2�.�W�������lW��1��D���1�0�&�y�w�}�W������F��Q1��D��
�
�
�0�{�}�W���Yӗ��X��B��*��e�0�d�$�{�}�W���YӇ��A��N��U���
�
�c�e�2�l��������9F�N��U���u�k�7�3�b�l�E߁�&¹��JǻN��U���0�u�k�7�1�h�F��&����D��=N��U���u�d�h�u�"��(��I����l��dךU��� �
�
�d���(���Y����\��CN��3���c�
�
������&����V9��N�����'�6�8�%��}�W���YӢ��R1��C��K��y�u�u�u�w�����
����VF�Z�U���u�u��1�2�.����Y���l�N�����4�u�_�u�w�}�W���Y����C9��\BךU���u�u�0�0�w�c����
��ƹF�N�����&�e�h�u�"��(��&����R��R��Y���u�u�u�6�g�`�W���&ƹ��9��1��E�ߊu�u�u�u�g�`�W���&ƹ��9��1��Y���u�u�u�4�3�8����Gӄ��lS��^��*ڊ�1�'�&�d�]�}�W���Y����X��B��*��
�
�
�0�{�}�W���Yӑ��[�U��@��e�0�e�"�f�W�W���Y�ƨ�[�U��@��e�0�e�1�~�W�W�������l_��h��*���u�:�%�;�9�}�6��I����lV��h[�� ���
�e�
�
�]�}�W�������^��d��U���u��!��3�5�J���K���F�N�����&�4�2�u�i�i�}���Y���r��R�����u�k�g�_�w�}�������9F�N��U���u�k�4�
�;�q�W���Y����V��S����&�y�u�u�w�}��������X��B��*��
�
�
�1�%�.�G�ԜY���F��N��U���
�
�d�
�����Y���F��N��U���
�
�d�
���G�ԜY���F��S�����k�7�3�`�n�m��������@��=N��U���u�0�u�k�5�;�B��I����l��d��U���u�"�d�h�w�(�(ځ�Hù��9��BךU���u�u�d�h�w�(�(ځ�Hù��9��UװU���7�3�`�d�d��(߁�Y�Ư�^��R �����a��c�
���(���&ƹ��9��d��Uʲ�;�'�6�8�'�u�W���Y����R��^
��U��f�y�u�u�w�}�6�������]��
P��Y���u�u�u��3�8�������T�N�����u�4�u�_�w�}�W��������T�����u�u�u�0�2�}�IϿ�&����9F�N��U���'�&�e�h�w�(�(ځ�J�Փ�lV��S
����_�u�u�u�w�8�W�������lW��1��E���e�_�u�u�w�}�G��Y����9��]��*ڊ�e�_�u�u�w�}����
���F��Q1��D��
�
�
�1�%�.�F�ԜY���F��N��U���
�
�f�f�2�m���s���F�@�H��� �
�
�f�d�8�G���H���F�N��U��7�3�`�d�d��(߁�H��ƓF�U��@��f�
�
�
�w�}��������^'��^��C���
�
�
� ���Gځ�&���F��Y��ʸ�%�}�u�u�w�}�3���.����[�\�U���u�u��1�2�.����Y���l�N��Uʔ�1�0�&�<�#�}�I��s���C	����U�ߊu�u�u�u�;�}�IϿ�&����9F�N��U���0�u�k�4��.�[���Y�����E��E��u� �
�
�d�n��������@��=N��U���u�0�u�k�5�;�B��J����9��BךU���u�u�e�h�w�(�(ځ�J�Փ�lW��BךU���u�u�1�'�$�l�J�������U��h��*���'�&�d�_�w�}�W��������h[��F���0�d�6�d�]�}�W���Y����X��B��*��f�0�d�"�f�W�W���Y�ƨ�[�U��@��f�
�
�
�f�f�}���Y����9��]��*؊�u�u�:�%�9�3�W���O�֊� ��h��*���
�
�e�
��W�W�������PF��GN��U���u�u��!� �9���Y����F�N��4���0�&�4�2�w�c�C�ԜY���F��S�����!�u�k�g�]�}�W���Ӌ��NǻN��U���9�u�k�4��1�[���Y�����R��Kʴ�
�&�y�u�w�}�WϿ�����F���*ߊ�f�f�0�g�6�9����U���F���U��7�3�`�d�d��(݁���ƹF�N��E��u� �
�
�d�n������ƹF�N�����&�d�h�u�"��(��J����l��E��D�ߊu�u�u�u�2�}�Iϼ��ӓ� U��R1����_�u�u�u�w�8�W�������lW��1��G���d�_�u�u�w�}�F��Y����9��]��*؊�d�n�_�u�w�)�B��A˹��	F��Z�����8��a��a��(���&����lW��d��Uʲ�;�'�6�8�'�u�W���Y����R��^
��U��f�y�u�u�w�}�6�������]��
P��Y���u�u�u��3�8�������T�N�����u�4�u�_�w�}�W��������T�����u�u�u�0�2�}�IϿ�&����9F�N��U���'�&�e�h�w�)�B��A˹��W��D^�U���u�u�6�e�j�}����H����P��=N��U���u�e�h�u�#�h�F��&����F�N�����0�&�u�k�;��(��A����A��BךU���u�u�0�u�i�1�(ځ�O�ޓ�VW�N��U���"�d�h�u�#�h�F��&����9F�N��U��h�u�!�`�f�e�(��s���F�F_��Kʹ�
�
�c�m�&�t�}���Yӊ��9��X��*ڊ�u�u�:�%�9�3�W���O�֊� ��h��*���`�d�m�_�w�}�����ơ�CF�N��U����!��1�?�`�W��s���F�v
�����4�2�u�k�c�W�W���Y�ƍ�W��D9�����k�g�_�u�w�2�ϳ�	��ƹF�N�����k�4�
�9�{�}�W���YӔ��V�	N��*���y�u�u�u�w�<����
���
��1�A܊�
�
�1�'�$�m�}���Y���P��
P�����d�a�
�
��8�[���Y�����
P�����d�a�
�
��m�}���Y���R��R��U��9�
�
�m�a�8�G�������JǻN��U���0�u�k�9���O����֓�VW�N��U���"�d�h�u�#�h�F��&����D��=N��U���u�d�h�u�#�h�F��&����WW�N��U���$�u�k�9���O����֓�O��=N��U���`�d�a�
���W�������V��Z/��Aړ�c�
�
�
��)�B��A���F��Y��ʸ�%�}�u�u�w�}�3���.����[�\�U���u�u��1�2�.����Y���l�N��Uʔ�1�0�&�<�#�}�I��s���C	����U�ߊu�u�u�u�;�}�IϿ�&����9F�N��U���0�u�k�4��.�[���Y�����E��E��u�!�`�d�c��(ށ�����@V�N��U���6�e�h�u�#�h�F��&����P��=N��U���u�e�h�u�#�h�F��&����BV�N��U���4�1�0�&�w�c����&����l��h�����d�_�u�u�w�}����Gӊ��9��X��*ۊ�0�y�u�u�w�}� ��D�Ơ�lS��Z�����"�d�_�u�w�}�W��D�Ơ�lS��Z�����1�y�u�u�w�}����Gӊ��9��X��*ۊ�d�n�_�u�w�)�B��@ƹ��9��N�����0�!�8��c��A���&����Q��1�@���e�u�u�2�9�/�ϳ�	��ƹF�N�����<�!�u�k�d�q�W���Y����W��D�����h�u�y�u�w�}�Wϟ�����d��_N��U���u�u�%�'�w�<�W�ԜY���F��\N��U���6�>�_�u�w�}�W��������E�����u�u�u�1�%�.�G��Y����lS��1��E���1�0�&�y�w�}�W������F��h[��C���0�e�6�e�]�}�W���Y���F��h[��C���0�e�$�y�w�}�W�������@��
P�����`�l�
�
��9����H���F�N��D��u�!�`�`�n��(߁���ƹF�N�����k�9�
�
�a�h��������F�N�����k�9�
�
�a�h��������9F���@���l�
�
�
�w�}��������^'��^��C���
�
�
� ���Gځ�&���F��Y��ʸ�%�}�u�u�w�}�3���.����[�\�U���u�u��1�2�.����Y���l�N��Uʔ�1�0�&�<�#�}�I��s���C	����U�ߊu�u�u�u�;�}�IϿ�&����9F�N��U���0�u�k�4��.�[���Y�����E��E��u�!�`�`�n��(ށ�����@V�N��U���6�e�h�u�#�h�B��&����P��=N��U���u�e�h�u�#�h�B��&����BV�N��U���4�1�0�&�w�c����&����l��h�����d�_�u�u�w�}����Gӊ��9��[��*ۊ�0�y�u�u�w�}� ��D�Ơ�lS��W�����"�d�_�u�w�}�W��D�Ơ�lS��W�����1�|�_�u�w�1�(ځ�O�ӓ�lT��T�����;�;�u��a�m�Fٸ�I����l��h[��Eߊ�
�_�u�u�2�8�������F�N��1����1�=�h�w�o�}���Y���r��R�����u�k�a�_�w�}�W�������@1��C��K��_�u�u�:�#�0����Y���F��[��Kʴ�
�9�y�u�w�}�WϬ�
���F��h��Y���u�u�u�4�3�8����Gӊ��9��[��*؊�1�'�&�e�]�}�W���Y����X��C1��@��
�
�
�0�{�}�W���Yӗ��X��C1��@��
�
�
�e�]�}�W���Y����V��S����
�c�`�0�e�<����
��ƹF�N�����k�9�
�
�a�h��������F�N����h�u�!�`�b�d�(���&����9F�N��U��h�u�!�`�b�d�(���&���9l�N�����d�m�
�u�w�2�����ơ�uP��q_��*ڊ�
�
� �
��e�C���YӁ��V����U�ߊu�u�u�u�6�<����Y���JǻN��U���1�'�&��9�8�J���U���F�/������1�=�h�w�t�W���	����^��d��U���u�6�>�h�w�-����s���F�E����u�%�'�!�]�}�W���Y����V��S����`�d�m�
�3�/���s���F�T�H��� �
�
�m�c�>�G�ԜY���F��S����`�d�m�
�g�W�W���Y�ƭ�W��D_��Kʷ�3�`�d�m��9����H���F�N��D��u� �
�
�o�i���s���F�@�H��� �
�
�m�c�*�F�ԜY���F��S����`�d�m�
�f�f�}���Y����U��Q��*���&�f�;�
�e�n����&����fW��N�����0�!�8��c��A���&����U��h]����;�
�g�f�1�1�(���s���T��E�����}�u�u�u�w��W���H���F�N��8�����h�u�{�}�W���Yӂ��9��s:��H���g�_�u�u�w�}����.����[�\�U���u�u�1� ���#���G����9F���ʸ�%�}�u�u�w�}����D�ƭ�l��d��U���u�'�&�!�j�}�������F�N�����k�2�%�3��h�B���U���F�
��D��u�'�
� �f�m�(��s���F�X�����k�2�%�3��h�B�������9F�N��U���h�u�'�
�"�l�Gځ����F�N�� ���k�2�%�3��h�B���P��ƹF��h^�����f�;�
�g�$�n�(ށ�����C9��N����:�0�!�8��i�1���&ù��F
�� ��Fػ�
�g�d�8�/�9����YӁ��V����U�ߊu�u�u�u��`�W��Y���F��b#��!���u�k�d�_�w�}�W����֓�z"��S�F���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���K���F��E�����_�u�u�u�w�4�G��Y����U��_�����u�u�u�u�3�3�W�������F9��Z��D�ߊu�u�u�u�8�)�J�������lW��1��\�ߠu�u�3�e�1�0�(���
����@9��1��E��6�8�:�0�#�0�1��?�Ъ�9��Z��G���f�;�
�
�]�}�W�������^��d��U���u��u�k�f�W�W���Y�Ƃ�~9��v)��H���y�u�u�u�w�9�߁�0����X�BךU���u�u�<�d� ��?��Y����F�N�����
���u�i�l�}���Y������FךU���u�u�<�e�j�}��������
9��d��U���u�1�;�u�i�:����&����l��=N��U���u�%�:�0�j�}��������
9��T��Y���u�u�u�1�"�}�IϹ�	����S��h�N�ߊu�u�
�
�4�-�Dݰ�&�Ԣ�lW��h;�U���:�%�;�;�w��A���Hŀ��l ��G1����g�&�d�d�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�t�W���	����^��d��U���u�1�;�u�i�;�(���<����G9��h��D��
�f�_�u�w�}�W���H���Q��1�Gڊ�
�
�e�_�w�}�W���	����[�C��F܊� �d�g�
�'�2��ԜY���F��B��Kʡ�%�f�
� �f�o�(��B���F��1�����g�&�f�;���(��Y�Ư�^��R �����a��c�
��>�������]��h_ךU���0�0�<�u�6�}�}���Y���z"�	N����u�u�u� ��	�0���G����F�N�����
���u�i�n�[���Y�����1��1���h�u�g�_�w�}�W�������z"��S�D�ߊu�u�:�!�:�-�_���Y�����N��U�������#�h�(���H����CU�N��U���1�;�u�k�5�;�B��Kù��9��d��U���u�:�6�1�w�c����M����lW��1�����y�u�u�u�w�9����GӒ��lR��Q��@���%�|�_�u�w�;�G�������]�� ��D��� �f�o�6�:�2�������� ��Q1�����
�g�&�f�9��(�ԜY�ƫ�]��TN�����u�u�u�u��}�I��s���F�y;��&����h�u�y�w�}�W�������d/��N��U��_�u�u�u�w�4�F���=���F��d��U���u�1� �
��	�W���H���F��E�����_�u�u�u�w�4�G��Y����v*��c!��*���3�
�c�c�'�q�W���Y����Z��
P�� ���
�c�e�0�f�,�[���Y���	��X
��H���8�
�b�3��h�B�������9F�N��U���!�h�u�8��j����L�ӓ�O��=dװ���u�x�!�0�4�/����
����N��h-�����u�3�!�0�$�<�ϳ�����F�=N��U����
�&�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����s���F�N��U���u�u�4�
��;���Y����`9��ZUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W������\��C��*��
�
�0�
�c�d�����Ƽ�\��D@��X���u�4�'�;�3�����K�ѓ�l��h_�L���&�2�
�'�4�g�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F�N��Uʴ�'�;�1�
�2�0�E�������lW��N�U���
�:�0�!�%��F؁�&¹��T9��_�U���u�u�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��@���!�0�u�u�w�}�W���Y���F���*���0�!�'�
�f��(���&����Z�V�����
�#�
�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C��D���2�d�c�u�$�4�Ϯ�����F�=N��U���'�2�d�c��.����	����	F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����	����l��h_�A���=�;�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��D���8�d�|�u�?�3�}���Y���F�N��U���<�
�0�
�c�l�K���	����@��A]��N���u�u�u�u�w�}�Wϻ�
���R��^	�����l�`�u�=�9�W�W���Y���F�N��Uʼ�
�0�
�a�f�a�W���&����_��G\�U���u�u�u�u�w�}������ƹF�N��U���;�u�3�u�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������T9��]�����;�%�:�0�$�}�Z���Yӏ��A��Z�*���<�;�%�:�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�e�|�!�2�}�W���Y���F�N��U���g�'�2�d�o�}�JϷ�J����lT��UךU���u�u�u�u�w�}����Y�έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���u�=�;�_�w�}�W���Y���F�N��*���
�a�f�i�w�-��������lV��N��U���u�u�u�u�2�9���Y���F�N�����3�u�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�܁�����
R��D��ʥ�:�0�&�u�z�}�WϷ�&����R��h�����%�:�u�u�%�>��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�r�p�}����Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W����έ�l��h��*��m�u�=�;�]�}�W���Y���F�N��ي�0�
�a�a�k�}��������ET��d��U���u�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*���� U��D��G���!�0�u�u�w�}�W���Y���F������d�l�u�h�>�i����K����9F�N��U���u�u�u�;�w�;�}���Y���F�R ����_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w���������\��h��*��g�4�&�2�w�/����W���F�^"�����'��:�
��8�(��K����Z��G��U���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���N����lT��N�����u�u�u�u�w�}�W���Y����9��h(��*���%�&�'�2�f�j�W������l ��h"����
�0�
�`�e�W�W���Y���F�N�����}�4�
�:�$�����&���R��^	������
�!�c�1�0�F���Y����l�N��U���u�u�u�u�w�4�(���?����\	��D1����b�u�h�4��2��������9F�N��U���u�u�u�;�w�;�}���Y���F�R ����_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�����M����@��YN�����&�u�x�u�w�4����H����R��P �����o�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��G�����_�u�u�u�w�}�W���Y���Z9��P1�F���h�<�d�'�0�o�A��Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���&����R��R�����:�&�
�#��f�W���Y���F�N�����3�_�u�u�w�}�W����ƥ�FǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���Ĺ��^9��G�����u�u�u�u�w�}�W�������\��C��*��
�
�
�0��i�F��Y����]	��h����b�<�d�3��h�@���B���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������A	��D�X�ߊu�u�'�6�$�}������ƹF��R	�����u�u�u�3��-���������������h�r�r�u�?�3�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�g�~�}����Y���F�N��U���9����#�/�(����ԓ�V�� Y�I���9����#�/�(����ԓ�F9��[��F�ߊu�u�u�u�w�}�W���*����^��R	��B��i�u�'�
�"�l�Fہ�K���F�N��U���u�3�
������&����Q��R�����3�
�`�`�'�f�W���Y���F�N��&��� ��;� ��i�F�������F�������;� �
�c�l����I�Փ� ]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��@���Y����9F�N��U���u�u�u�9���/�������S��R1�����g�g�u�h�;��(��O����l��=N��U���u�u�u�u�w�1�>���!����V��[�����'�2�g�f�w�`����&����l��h����u�u�u�u�w�}�W���0����r4��R��D���0�e�'�2�e�n�W������^��h��*��_�u�u�u�w�}�W���Y����}"��v<�����d�g�0�d�%�:�E��Y����G9��V�*���
�d�_�u�w�}�W���Y���U5��y*��4���0�8�b�
�2��O��E�Ơ�lS��V����u�u�u�u�w�}�W�������w#��e<�����b�'�2�g�f�}�Jϲ�&ƹ��^��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�e�����A���G��=N��U���u�u�u�u�w�1�>���!����V��[�����'�2�g�b�w�`����&����l��h����u�u�u�u�w�}�W���0����r4��R��D���0�d�'�2�e�e�W������^��h��*��_�u�u�u�w�}�W���Y����}"��v<�����d�c�0�e�%�:�E��Y����G9��V�*���
�d�_�u�w�}�W���Y���P
��y*��4���0�8�d�c�2�l����K����[��C1��D��
�
�
�d�]�}�W���Y���F�Q=��;�����0�8�`�����A���F��h[��C���$�n�u�u�w�}�W���Y����`9��s+��'���'�
�d�'�0�o�@���Dӊ��9��V��D�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Eځ�
����O�C�����u�u�u�u�w�}�W�������A9��X��F���e�'�2�g�n�}�Jϼ��ӓ� U��R1����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C�����;�%�:�0�$�}�Z���YӖ��P��F��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y�����Yd��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O������u�u�u�u�w�}�WϽ�&����\��X��Gي�
�
�0�
�a�n�K�������U��h��*��_�u�u�u�w�}�W���Y����G9��E1�����l�0�e�'�0�o�N���Dӄ��lS��\�����$�n�u�u�w�}�W���Y����_9��h(��*���%�g�
�
��8�(��L���Q��1�Gڊ�
�
�e�_�w�}�W���Y���F��h=��0��� �
�c�'�0�o�F���DӀ��`#��t:�����
� �d�g��n�}���Y���F�N�����!�%�d�<�%�:�E��Y����V
��Z�*��� �d�a�
�e�W�W���Y���F�N�����%�e�<�'�0�o�D���Dӕ��l��^��*���d�b�
�g�]�}�W���Y���F�D�����l�<�'�2�e�i�W��
����^��h�� ��m�
�g�_�w�}�W���Y���F��[1�����<�'�2�g�c�}�Jϭ����� Q��h��D��
�g�_�u�w�}�W���Y���G��\�����b�m�i�u�:��E���&����l��=N��U���u�u�u�u�w�0�(�������T��S�����m�3�
�m�b�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�|�u�?�3�W���Y���F�N��&��� ���!��1����&�ԓ�V�� V�I���'�
� �d�f��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��E���8�d�|�|�#�8�}���Y���F�N��������!�b�����O���F��G1��*���`�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���=�;�u�u�w�}�W���Y����9��h(��*���%�d�
�0��h�E��Y����Z9��E1�����m�3�
�c�c�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����d�|�u�=�9�}�W���Y���F���*���
�a�d�i�w��(���H����CT��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�e�1�0�E���PӒ��]l�N��U���u�u�u�<�d�/���@�����h��G��
�g�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��_��\ʡ�0�_�u�u�w�}�W���Y�ƥ�9��P1�G���h�<�a�3��o�D���B���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������A	��D�X�ߊu�u�'�6�$�}������ƹF��R	�����u�u�u�3��-���������������h�r�r�u�?�3�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�d�g�`��������l��R	��B��u�;�u�4��2����¹��F��[1�����<�'�2�g�d�t����Q����\��h��*���u�0�
�8�e��(���&����F��SN�����;�!�9�d�g�`��������l��R	��B��u�;�u�4��2��������F�V�����&�$��
�#�k����K�����Yd��U���u�u�u�u�w�-����&����T9��^��Hʥ�<�8�
�
�"�o�Bׁ�J���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���b�3�8�d�~�<����	����@��A_��U���-�!�:�1��(�F��&���F��R ךU���u�u�u�u�w�}�W�������l��h\�B��1�"�!�u�~�a�W���&�Փ�F9��^��D��1�"�!�u�~�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�4�1�}�'�>�����ד�[��R����
�
�0�
�`�d�W���Yۇ��P	��C1��D��h�&�9�!�'�m��������O��Y
�����:�&�
�#��}�W���&����
9��E��G��|�4�1�}�'�>�����ד�[��R����
�
�0�
�`�j�W���Yۇ��P	��C1��D��h�!�%�a��8�(��J���G��=N��U���u�u�u�u�w�0�(�������P��S�����b�3�
�d�d�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�l�u�;�w�<�(���
����9��
N�����;�d�3�
�f�e����PӒ��]l�N��U���u�u�u�u�w�)���&����_��\�����:�e�u�h�#�-�C߁�����9��\�����:�e�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h]�U���u�4�
�:�$��ށ�Y�Ʃ�Z��Y
�� ��e�
�g�|�w�5����Y���F�N��U���u�8�
�d�%�:�E��Q�ƨ�D��^��I���8�
�d�3��o�N���Q�ƨ�D��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o����H�ƭ�WF��O�����
� �d�a��o�JϿ�&����G9��1�\���=�;�u�u�w�}�W���Y���F��Z�����a�c�g�1� �)�W���E�Ƹ�C9��h_�A���}�u�:�;�8�m�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u� ���Bց�����V��]�Dʱ�"�!�u�|�k�}�G���s���Q��1�Cӊ�1�'�'�2�e�i�_�������V�S��E���_�u�u�!�b�l�Oׁ�����V��Z�Dʱ�"�!�u�|�k�}�G���s���Q��1�Mފ�1�'�'�2�e�h�_���E���]ǻN�����0�
�a�c�a�}�������[�^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����l�N����
�0�
�`�`�k�W������F�L�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����D��N�����a�
�0�
�n�i�A�������U�S��E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��d��Uʡ�%�a�
�0��d�C��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�����u�x�u�=�w�8�ϭ����R��d1�����3�!�0�&�6�8�������KǻN�����
�&�
�&�>�3����Y�Ƽ�\��DN�����4�!�u�%���������F��h�����
�0�1�'�6����M������C��ߊ� �d�a�
�e�}��������U��X�����0�<�6�;�d�;�(��@������C��؊� �d�e�
�e�}��������U��V�����0�<�6�;��(�E��&���F�U�����u�u�u�6�$�}����&����ZǻN��U���u�u�=�;�6��#���H����lV�	NךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ��έ�l��E��U���6�;�!�9�0�>�G���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=�����3�8�d�_�w�}�W���Y���F��DךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����3�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]°�<�6�;�`�1��B���	���R��X ��*���
�|�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����l ��h]�U���u�u�u�u�w�}�������R��X ��*���<�
�u�u�'�>�^Ͽ��Ω�Z��Y
�����`�g�%�u�w�-��������lV�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!��.�(��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�E�������F�N��U���u�u�0�1�>�f�W���Y���F��_������&�f�3�:�o�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���J����lT��N��U���u�u�u�u�2�9���Y���F�N�����4�
��&�c�;���D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����l ��h]�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�B������FǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���O����lS�	NךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��C�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����]��QUךU���u�u�u�u�?�3����-����l ��hX��K�ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��h�����#�
�u�u�/�)����&����P��G\��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�N�������F�N��U���u�u�0�&�1�u�_�������l
��^��U���%�6�|�4�3�u��������EW��S�����:�1�
� �f�k�(��P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��[��U���u�u�u�u�w�}�W�������l ��R������&�b�3�:�k�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��M���8�b�h�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�o�;���s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���l�3�8�m�j�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�g�;���s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���ց�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�e�1�0�N��Y���F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��D��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��Dۊ�&�
�e�_�w�}�W���Y���F��SN��N���u�u�u�u�w�*����	����@��h��*��h�u�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����&�!�e�'�6���������9��S�����;�!�9�d�g�t����Q����\��h��*���u�-�!�:�3����Aʹ��O�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�g�1�0�F��Y���F�N��U���9�<�u�}�6�����&����P9��
N��*���u�;�u�}�9�/����I����W9��V
�� ��a�%�u�u�'�>�����ד�F�� ��]´�
�:�&�
�!��W�������]��Q��@���%�|�|�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����U��D��G�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��G���8�d�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GW��Q��D���k�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�f�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�f�1�0�F��Y���F�N��U���;�u�3�_�w�}�W���Y�ƻ�V��G1��*���a�3�8�d�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�����M���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���M����lW��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�h����H���l�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��[�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��[�����a�_�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�"�2�}����&����l ��h_�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��B���8�d�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�d�
�&��h�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��D݊�&�
�c�h�w�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�%�6�;�#�1�F��DӃ��G��S\�� ��e�
�g�|�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�d�e�h�2�4����K����P��h�\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Fׁ�
����l�N��U���u�u�u�0�$�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����l ��h_����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��D��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��DҊ�&�
�b�_�w�}�W���Y���F��SN��N���u�u�u�u�w�*����	����@��h��*��h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���e�3�8�d�l�}�W���Y���F������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d��.�(��s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���g�
�&�
�n�`�W���Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�l����K��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���Kù��^9��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���;�4�
��$�o�(���&���FǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����l ��h\����u�u�u�u�w�}�W������F�N��U���u�u�u�%������DӇ��`2��C\�����g�n�u�u�w�}�W���Y����]��QUךU���u�u�u�u�?�3����-����9��Z1�U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��Gي�&�
�g�_�w�}�W���Y���F��DךU���u�u�u�u�w�}�W���	����U��S�����
�!�g�3�:�o�L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:�����3�8�g�u�i�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�g��.�(��s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!�c�;���Y���F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���Kƹ��^9��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$����ӓ�@��N��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�%������DӇ��`2��C\�����g�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���g�
�&�
�c�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�`�h�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�b�3�:�o�L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�o�(���&����F�N��U���u�u�0�1�>�f�W���Y���F��_������&�g�
�$��A��Y���F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	���&����Q�	NךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�g�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��1����u�k�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����*����Z�V��!���f�
�&�
�n�W�W���Y���F�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�n�;���B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�e�3�8�e�}�I�ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�4��2����¹��F��^�����3�
�d�m�'�t�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��G���8�f�n�u�w�}�W���Y�����^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�#��}�W�������9��h\�M���|�|�!�0�]�}�W���Y���F�N������3�8�i�w�-�$����ד�@��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�=�9�<�(���
����U��^��K�ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�4������E�ƭ�l5��D�*���
�l�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�d�3�8�d�f�W���Y���F�N�����3�_�u�u�w�}�W�������C9��h��G���8�f�u�k�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����4�
�:�&��+�(���Y����P	��h��G��
�g�|�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����e�h�0�<�4�3�(���K����CT�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�d�;���B���F�N��U���u�9�0�u�w�}�W���Y���F���;���&�u�h�4��	���&���� W��N��U���u�u�u�u�2�9���Y���F�N�����4�
��&�d�����K���9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N������3�8�i�w�-�$����ԓ�@��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�=�9�2����Y���9F�N��U���u�u�u�%������D�Ĕ�k>��o6��-���������/���!���9F�N��U���u�4�0�_�w�}��������@]ǑN��X���%�1�;�u�$�4�Ϯ�����F�=N��U���1�;�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1�U���6�y�4�
�>�����*���� T��D��D���-�!�:�1�1��E���	��ƹF��R	�����u�u�u�3��u��������]��[����h�4�
�!�%�t�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�f�
�$��F����Ƣ�GN��G1�����9�d�e�h�2�4����&����V��G\��\���!�0�u�u�w�}�W���YӇ��W	��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�9����DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W�������R��P �����&�{�x�_�w�}��������@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�W�W�������F�N�����}�:�}�4��2��������F�V�����|�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&�����YNךU���u�u�u�u�'�4����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����1�0�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�0�3�}����Ӗ��P��N����u�%�'�4�.�<����&����\��E�����%�6�y�4��4�(�������@��h��*��u�-�!�:�3�;�(��N����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&���� W�V �����}�%�6�;�#�1�F��DӃ��G��S1��*��b�%�|�|�w�5��ԜY���F�N��*���1�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����V��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����C9��C��*���h�6�
����%�������l��h��*��c�_�u�u�'�/����&�����~ ��-���!�'�
�`���(���&����l�N��*��� �;�d�u�j�;�(���<����G��hY�����g�c�n�u�w�<�(�������F���<�����!�'��l����K����9F������'�
�u�h�4��9���8����A��\��*ڊ�0�
�m�c�]�}�W�������]9��S��������!�%��B݁�&¹��T9��_�U���4�
�0� �9�i�K�������v>��e����a�0�e�'�0�o�@��Y����C9��C��*���h�6�
����%�������l��h��*��d�_�u�u�'�/����&�����~ ��-���!�'�
�`���(���&����l�N��*��� �;�b�i�w�1�>���!����V��[�����'�2�g�l�l�}�WϿ�&����A��R���������2�0�@؁�����W��N�����0� �;�l�k�}�$���=����a��Z1�*���
�m�`�_�w�}�Z���	����l��h_�U���<�;�%�:�2�.�W��Y����C9��P1����f�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����f�i�u�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��CF�����4�!�h�4��2��������O�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����l�u�&�<�9�-����
���9F������7�1�d�l��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��N�����T�����d�d�h�4������H�ƨ�D��_�\�ߊu�u�;�u�%�>���s���K�V�����1�
�l�a�6�.��������@H�d��Uʴ�
�<�
�1��d�C���
����C��T�����&�}�%�6�{�4�(�������A��h�����
�l�
�g�]�}�W������F�N��U���u�4�
�<��9�(��M���N��h�����:�<�
�u�w�-��������\�^ �����
�
�0�1�%�<�(���K�ғ�F�V�����
�#�
�|�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����@����@��YN�����&�u�x�u�w�<�(���&����_��h�����%�:�u�u�%�>����	����l��F1��*���g�3�8�d�{�8�����Փ�F9��W��G�ߊu�u�0�<�]�}�W���Y���F�V�����1�
�l�`�k�}�_�������l
��^��U���%�&�2�6�2��#���H����^9��N�����%�6�;�!�;�l�G������\��h��D��
�g�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��N������]F��X�����x�u�u�4��4�(���&����l��^	�����u�u�'�6�$�u��������B9��h��E���8�g�y�0�>�>��������^��GךU���0�<�_�u�w�}�W���Y���R��^	�����l�m�i�u��-��������Z��S�����2�6�0�
��.�D߁�
����F��SN�����%�6�;�!�;�l�G������\��h��G��
�g�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��]�I���4�
�:�&��+�(���Y����`9��ZF����!�u�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��[�I���4�
�:�&��+�(���Y����`9��ZF����!�u�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��X�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�d�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���HӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�D��u�4�
�:�$��ށ�Y�ƭ�l%��Q��D���:�;�:�d�~�f�W�������A	��D����u�x�u�%�$�:����J����@��YN�����&�u�x�u�w�<�(���&���� V��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��F���i�u�4�
�8�.�(���&���R��d1����u�:�;�:�f�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����l�i�u�4��2����¹��F��h-�����d�u�:�;�8�l�^��Y����]��E����_�u�u�x�w�-�������� U��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��]�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����f�f�i�u�6�����&����F�V��&���8�d�u�:�9�2�F���B����������n�_�u�u�z�}��������lU�������%�:�0�&�w�p�W�������T9��S1�A���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�a�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W�� X�����;�%�:�0�$�}�Z���YӇ��@��U
��F���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�f�c�k�}��������_��N������3�8�d�w�2����H���9F���U���6�&�n�_�w�}�Z���	����l��h]�U���<�;�%�:�2�.�W��Y����C9��P1����m�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�f�o�a�Wǿ�&����G9��1�Hʴ�
��3�8�e�}��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��E���&�<�;�%�8�8����T�����D�����a�m�4�&�0�����CӖ��P����6���&�|�u�u�5�:����Y���F�N��U���&�2�7�1�c�e�K�������]��[��D��4�
��3�:�o�W������O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�a�l�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�i�N��Yۇ��P	��C1��D��h�4�
��1�0�E�������T��UךU���;�u�'�6�$�f�}���Y���R��^	�����c�u�&�<�9�-����
���9F������7�1�a�b�6�.���������T��]����
�&�|�w�}�������F�N��U���u�%�&�2�5�9�C��E����C9��Y�����d�h�4�
��;���Y����G	�G����u�;�u�'�4�.�L�ԶY���F��h��*���
�b�u�&�>�3�������KǻN�����2�7�1�a�o�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���A�����T�����d�d�h�4������K�ƨ�D��\�\�ߊu�u�;�u�%�>���s���K�V�����1�
�m�u�$�4�Ϯ�����F�=N��U���&�2�7�1�c�e��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����M���F��G1�����9�d�d�h�6��$�������W	��C��@���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�l�w�.����	����@�CךU���%�&�2�7�3�i�N���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(������F��@ ��U��|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�f�<����Y����V��C�U���4�
�<�
�3��F���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������[�V��&���8�e�1�"�#�}�^������]��[��D��u�u�0�1�'�2����s���F������7�1�`�e�6�.��������@H�d��Uʴ�
�<�
�1��n�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&����[�V�����
�#�
�u�w�-�4���
������Y��G���n�u�u�0�3�-����
��ƓF�C�����2�7�1�`�b�<����Y����V��C�U���4�
�<�
�3��Cځ�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&����_��X����|�n�u�u�2�9��������9l�N�U���&�2�7�1�b�k�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����P��S�����:�&�
�#��}�W���:����^N��
�����f�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�e�NϿ�
����C��R��U���u�u�4�
�>�����Iʹ��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��N�����u�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�e�GϿ�
����C��R��U���u�u�4�
�>�����Kù��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��N�����u�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�e�OϿ�
����C��R��U���u�u�4�
�>�����K˹��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U�� N�����u�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�e�GϿ�
����C��R��U���u�u�4�
�>�����Mù��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��^�����:�d�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�O������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��[�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�d�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@Ӈ��Z��G�����u�x�u�u�6���������
9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�4�
�:�$��ށ�Y�ƭ�l%��Q��G���:�;�:�g�~�f�W�������A	��D����u�x�u�%�$�:����A����@��YN�����&�u�x�u�w�<�(���&����P��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��M��i�u�4�
�8�.�(���&���R��d1����u�:�;�:�d�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����l�i�u�4��2����¹��F��h-�����f�u�:�;�8�n�^��Y����]��E����_�u�u�x�w�-��������
P��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��W�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����m�c�i�u�6�����&����F�V��&���8�f�1�"�#�}�^��Y����]��E����_�u�u�x�w�-��������P��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��^�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����l�c�i�u�6�����&����F�V��&���8�a�1�"�#�}�^��Y����]��E����_�u�u�x�w�-��������^��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��\�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����l�m�i�u�6�����&����F�V��&���8�m�1�"�#�}�^��Y����]��E����_�u�u�x�w�-��������W��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��Z�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����l�d�i�u�6�����&����F�V��&���8�l�1�"�#�}�^��Y����]��E����_�u�u�x�w�-��������`2��C_�����l�4�&�2�w�/����W���F�V�����&�$��
�#�m����@����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�l�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�d�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��D���8�d�u�&�>�3�������KǻN�����2�6�0�
��.�Fށ�
����l��^	�����u�u�'�6�$�u��������l^��d��Uʷ�2�;�u�u�w�}��������T9��S1�E���=�;�_�u�w�}�W���Y����Z��D��&���!�d�3�8�f�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�l����H�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�g�3�8�f�}����Ӗ��P��N����u�%�&�2�4�8�(���
����U��_�����;�%�:�u�w�/����Q����Z��S
��C���u�u�7�2�9�}�W���Yӏ����D�����g�b�u�=�9�W�W���Y���F��h��*���$��
�!�e�;���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���K����lW��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!�d�;���Y����T��E�����x�_�u�u�'�.��������l��1����
�&�<�;�'�2�W�������@N��h��*���
�l�|�u�w�?����Y���F��QN�����2�7�1�g�f�}����s���F�N�����<�
�&�$����������F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����U��D��G��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���������� F��D��U���6�&�{�x�]�}�W���
����@��d:�����3�8�d�
�$�4��������C��R�����<�
�1�
�g�t�W�������9F�N��U���}�%�&�2�5�9�D��Y����l�N��U���u�4�
�<��.����&����l ��h_�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(���&����l5��D�*���
�f�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��.����&����l ��h_����2�u�'�6�$�s�Z�ԜY�ƭ�l��h�����
�!�`�3�:�l�(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��[�����a�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���d�
�&�
�c�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9��X�����`�4�&�2�w�/����W���F�V�����&�$��
�#�k����Hƹ��@��h����%�:�0�&�6���������OǻN�����_�u�u�u�w�;�_���
����W��_�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�`�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�d��.�(��E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�c�6�.��������@H�d��Uʴ�
�<�
�&�&��(���N����lW��V�����'�6�o�%�8�8�ǿ�&����Q��]����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�d�
�$��A��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�F؁�
����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�d�
�$��@Ͽ�
����C��R��U���u�u�4�
�>�����*����^��D��B���&�2�
�'�4�g��������C9��P1����a�_�u�u�2�4�}���Y���Z �V�����1�
�c�|�#�8�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
����U��Y��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�l�(���&����@��YN�����&�u�x�u�w�<�(���&����l5��D�*���
�m�4�&�0�����CӖ��P�������7�1�d�l�~�}�Wϼ���ƹF�N�����%�&�2�7�3�l�N�������9F�N��U���u�%�&�2�4�8�(���
����U��V��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
�ד�@�������%�:�0�&�w�p�W�������T9��R��!���d�3�8�e�6�.���������T��]���&�2�7�1�b�t�W�������9F�N��U���}�%�&�2�5�9�B�������9F�N��U���u�%�&�2�4�8�(���
�ד�@��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	���&����_��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=����
�&�
�l�6�.���������T��]���&�2�7�1�d�k�}���Y����]l�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��E���8�d�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����9��Z1�U���<�;�%�:�2�.�W��Y����C9��P1������&�g�
�$��G���
����C��T�����&�}�%�&�0�?���A���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��C\�����g�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�d�3�8�e�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C\�����g�u�&�<�9�-����
���9F������6�0�
��$�o�(���&�ד�@��Y1�����u�'�6�&��-��������^�N�����;�u�u�u�w�4�Wǿ�&����Q��^�U���;�_�u�u�w�}�W���	����l��F1��*���g�3�8�g�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!�e�;���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���f�3�8�g�w�.����	����@�CךU���%�&�2�6�2��#���K����^9��h�����%�:�u�u�%�>����	����l��hZ�\���u�7�2�;�w�}�W�������C9��P1����l�u�=�;�]�}�W���Y���R��^	������
�!�f�1�0�E���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$����������F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�a�1�0�E���
������T��[���_�u�u�%�$�:����&����GT��Q��Gي�&�<�;�%�8�}�W�������R��^	�����c�|�u�u�5�:����Y����������7�1�a�b�w�5��ԜY���F�N��*���
�&�$���)�C�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����l ��h\�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�B�������R��P �����&�{�x�_�w�}��������B9��h��@���8�g�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�b�~�}�Wϼ���ƹF�N�����%�&�2�7�3�i�O������F�N��U���4�
�<�
�$�,�$����ӓ�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��[�����a�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����Г�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�c�3�8�e���������PF��G�����4�
�<�
�3��O���Y����V��=N��U���u�3�}�%�$�:����M���G��d��U���u�u�u�4��4�(�������@��h��*���i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�`�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*��4�&�2�u�%�>���T���F��h��*���$��
�!�`�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������l^��N�����u�u�u�u�w�}��������V��c1��G݊�&�
�c�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�g�
�$��A��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��GҊ�&�
�b�4�$�:�W�������K��N�����<�
�&�$����������9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��L���!�0�u�u�w�}�W���YӇ��@��T��*���&�g�
�&��j�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�o�(���&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�g�
�&��e�����Ƽ�\��D@��X���u�4�
�<��.����&����l ��h\�����2�
�'�6�m�-����
ۇ��@��U
��@��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�f�|�!�2�}�W���Y���F��G1�����0�
��&�e�����A���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���Kʹ��^9��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�e�;�������]F��X�����x�u�u�4��4�(�������@��Q��D���&�2�
�'�4�g��������C9��P1����e�_�u�u�2�4�}���Y���Z �V�����1�
�f�|�#�8�W���Y���F������6�0�
��$�o����H���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���K����lW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�f��.�(������]F��X�����x�u�u�4��4�(�������@��h��*���4�&�2�
�%�>�MϮ�������D�����`�`�_�u�w�8��ԜY���F��F��*���
�1�
�a�~�)����Y���F�N�����2�6�0�
��.�D߁�
����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�Dށ�
������^	�����0�&�u�x�w�}��������V��c1��Fۊ�&�
�e�4�$�:�(�������A	��D�����2�7�1�m�n�W�W�������F�N�����4�
�<�
�3��A�������9F�N��U���u�%�&�2�4�8�(���
����U��^��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C]�����f�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��_�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�f�
�&��l��������\������}�%�&�2�5�9�B��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���g�3�8�f�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�d�����K����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�f�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�f�1�0�D���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ي�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�D����ԓ�@��Y1�����u�'�6�&��-��������_�N�����;�u�u�u�w�4�Wǿ�&����Q��^�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��*���
�u�&�<�9�-����
���9F������6�0�
��$�i����J����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:��ފ�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C[�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�b�;��������]9��X��U���6�&�}�%�$�:����@���F�U�����u�u�u�<�w�<�(���&����
V�����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��h��*���&�<�;�%�8�8����T�����D�����
��&�c�1�0�B���
����C��T�����&�}�%�&�0�?���I���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��CX�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GQ��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�b�3�:�k��������\������}�%�&�2�5�9�E��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:��݊�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����l ��hY�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�m�3�8�`�<����&����\��E�����%�&�2�7�3�e�O�ԜY�Ʈ�T��N��U���<�u�4�
�>�����K����[��=N��U���u�u�u�%�$�:����&����G^��D��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
�ߓ�@�������%�:�0�&�w�p�W�������T9��R��!���l�3�8�m�6�.���������T��]���&�2�7�1�n�e�}���Y����]l�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�%�&�0�>����-����l ��hV��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��CW�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN�����:�0�!�'��l�(���&����P��G\��Hʦ�1�9�2�6�!�>��������V��E�����!�'�
�d������M���F��D�����%�6�;�!�;�o�F���s���Q��1�Fي�
�
�1�'�$�m�K�������l��h\�B��x�d�1�"�#�}�^�ԶY���F��Q1��D��
�
�
�1�%�.�FϿ�
����C��R��U���u�u�7�3�b�l�D܁�&ù��W��D_�����;�%�:�u�w�/����Q����Z��D��&���!�f�3�8�f�q��������V��c1��Dފ�&�
�f�u�'�.��������l��1����y�4�
�<��.����&����l ��h_����u�0�<�_�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*���|�!�0�u�w�}�W���Y����F ��h_�F���e�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�c�t����Y���F�N��U���
�
�f�f�2�m��������[��G1�����9�c�
�}�w�}�W������]ǻN��U���9�<�u�}�'�>��������lW������6�0�
��$�l�(���&�����YNךU���u�u�u�u�"��(��J����l��E��D��u�%�6�;�#�1�Aہ�Q���F��@ ��U���_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-���� 9��Z1�\���=�;�_�u�w�}�W���Y����9��]��*ڊ�1�'�&�d�k�}��������EP��F�X��1�"�!�u�~�W�W���Y�Ʃ�@�N��U���u�u�7�3�b�l�D܁�&ù��W��D_��H����n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϼ��ӓ� U��R1����4�&�2�u�%�>���T���F��Q1��D��
�
�
�0��.����	����	F��X��´�
�0�u�%�$�:����&����GT��Q��G���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��Z�����f�|�u�=�9�W�W���Y���F��Q1��D��
�
�
�0�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��Q1��D��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��J����l�������%�:�0�&�w�p�W�������lW��1��E���d�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���J����lW�������6�0�
��$�l�(���&���R��^	������
�!�`�1�0�F������T9��R��!���d�
�&�
�b�W�W�������F�N�����}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��E������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�'�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�b�;���P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��X�����`�|�|�!�2�}�W���Y���F��B��*��f�0�e�6�f�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��f�0�e�6�f�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�7�3�b�l�D܁�&ù��Z�U��@��`�0�e�$�l�W�W���Tӄ��lS��]�����"�d�4�&�0�}����
���l�N�����d�f�
�
��8�(�������A	��N�����&�4�
�0�w�-��������`2��C_�����d�y�4�
�>�����*����R��D��F���%�&�2�6�2��#���Hƹ��^9��N��*���
�&�$���)�A�������9F����ߊu�u�u�u�1�u�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���J����lW��N��U���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��Z��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�c�3�:�l�^���Y����l�N��U���u�7�3�`�f�n�(���&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�7�3�`�f�n�(���&����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W�������U��h��*���'�&�e�i�w�0�(�������Q��N�Dʱ�"�!�u�|�]�}�W��Y����9��]��*ۊ�1�'�&�d�6�.��������@H�d��Uʷ�3�`�d�f���(�������l��^	�����u�u�'�6�$�u��������B9��h��F���8�d�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
����U��Z����<�
�&�$����������OǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����Г�@��G�����u�u�u�u�w�}�Wϼ��ӓ� U��R1�����0�&�u�h�6�����&����lU�C��U���;�:�e�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�a�|�!�2�}�W���Y���F��B��*��f�0�d�4�3�8����DӇ��P	��C1��Cފ�}�u�u�u�8�3���B���F������}�%�6�;�#�1����H����C9��P1������&�d�
�$��D�������9F�N��U���u� �
�
�d�n��������@��S�����;�!�9�c��u�W���Y����G	�UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����T����ߊu�u�u�u�w�}����&����l��h�����d�i�u�%�4�3����Oǹ��F�N�����u�|�_�u�w�}�W������F�N��Uʷ�3�`�d�f���(�������Z�6��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�5�;�B��J����9��N�����u�'�6�&�y�p�}���Y����9��]��*ۊ�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���Kù��^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���=�;�_�u�w�}�W���Y����9��]��*ۊ�0�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����9��]��*ۊ�0�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u� �
�
�d�n��������@��YN�����&�u�x�u�w�?����H����V9��T�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�n����H����C9��P1������&�d�
�$��D���	����l��F1��*���`�3�8�d�{�<�(���&����l5��D�*���
�`�_�u�w�8��ԜY���F��F��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�g�~�2�W���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���Hǹ��^9��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�`�3�8�f�t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���!�0�u�u�w�}�W���Yӄ��lS��]�����6�d�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���Yӄ��lS��]�����6�d�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʷ�3�`�d�f���(��E�Ʈ�U9��^�����$�n�_�u�w�p����L���� 9��1��Dʴ�&�2�u�'�4�.�Y��s���Q��1�Fي�
�
�0�
�$�4��������C��R�����0�u�%�&�0�>����-���� 9��Z1�Yʴ�
�<�
�&�&��(���M����lW�������6�0�
��$�l�(���&���R��^	������
�!�c�1�0�F���Y����V��=N��U���u�3�}�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�n����H���\������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�|�:�w�u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fځ�
����O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�~�}����s���F�N�����`�d�f�
������DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����`�d�f�
������DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�(�(ځ�J�Փ�lT��S
����i�u�8�
�d�/���N����F��S�����|�_�u�u�z�}����&����l��h�����d�4�&�2�w�/����W���F�U��@��f�
�
�
�3�/��������]9��X��U���6�&�}�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����ғ�@��B�����2�6�0�
��.�Fځ�
����F��h��*���$��
�!�a�;���P�����^ ךU���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�A�������F��R ��U���u�u�u�u�5�;�B��J����9��S�����h�4�
�:�$�����J���W��X����n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����S��D��A���!�0�u�u�w�}�W���Yӄ��lS��]�����4�1�0�&�w�`��������_��h\��U���u�:�;�:�g�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�f�~�)����Y���F�N�� ���
�f�f�0�e�<����
�����T�����c�
�}�u�w�}�������9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����K����[��=N��U���u�u�u� ���D����ԓ�W��D�I���%�6�;�!�;�k�(���Y����W	��C��\�ߊu�u�u�u�;�8�}���Y���F�U��@��f�
�
�
�3�/���E����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�7�3�`�f�n�(���&����R��P �����&�{�x�_�w�}����&����l��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�o�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O����ߊu�u�u�u�w�}����&����l��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}����&����l��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�� ���
�f�f�0�e�>�FϿ�
����C��R��U���u�u�7�3�b�l�D܁�&����9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�f�3�:�l�[Ͽ�&����P��h=����
�&�
�f�w�-��������`2��C_�����d�y�4�
�>�����*����P��D��@�ߊu�u�0�<�]�}�W���Y���N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��]�����g�|�:�u��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��@���8�d�|�u�%�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O�N�����u�u�u�u�w�}����L���� 9��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����L���� 9��1��D��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�U��@��f�
�
�
�f�a�W���&ƹ��9��1��N�ߊu�u�x�7�1�h�F��&����D��V�����'�6�&�{�z�W�W�������U��h��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����T�V�����&�$��
�#�i����H����C9��P1������&�d�
�$��C���	����l��F1��*���c�3�8�d�~�}�Wϼ���ƹF�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�f�3�:�l�^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����R��D��F���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��PӉ��N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�|�u�=�9�W�W���Y���F��Q1��D��
�
�
�0�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��Q1��D��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u� �
��h�N�������C9��hZ�*��i�u�%�6�9�)���&����F��S�����|�_�u�u�"��(��@����A��N�U���
�f�3�
�a�m����Y����W	��C��\�ߠu�u�x�u�"��(��@����A��N�����u�'�6�&�y�p�}���Y����9��W�����&�d�4�&�0�����CӖ��P����*ߊ�`�l�4�1��8�(��J�ƭ�l��h�����
�!�
�&��q��������V��c1��M���8�b�u�%�$�:����&����GR��D��Yʡ�%�g�
� �f�e�(��s���Q��Yd��U���u�<�u�}�'�>��������lW������6�0�
��$�e����N����[��=N��U���u�u�u� ���B�������@��S�����d�3�
�`�c�-�_���Y�ƨ�D��^����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���M����lU����ߊu�u�u�u�w�}����&����l��E��D��u�%�6�;�#�1�Aہ�Q���F��@ ��U���_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����l ��h_��U���;�_�u�u�w�}�W�������S��h�����d�i�u� ���B�������A��Z�N���u�u�u�0�$�}�W���Y���F��B��*���l�4�1�0�$�}�J���!��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�`�l�4�m�����Ƽ�\��D@��X���u�7�3�`�f�k�(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�d�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�a�t�W������F�N��Uʷ�3�`�d�c��8�W������]��[����_�u�u�u�w�1��ԜY���F�N�����d�c�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��@������^	�����0�&�u�x�w�}����L����
9��1�����
�'�6�o�'�2��������F��h��*���$��
�!��.�(������T9��R��!���m�3�8�b�w�-��������`2��CZ�����|�u�u�7�0�3�W���Y����UF�F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&���\������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����f�|�|�!�2�}�W���Y���F��B��*���l�6�d�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����F ��h_�L���d�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���7�3�`�d�a��FϿ�
����C��R��U���u�u�7�3�b�l�Aց�H����Z��G��U���'�6�&�}�9��(ށ�&����]9��h_��*���3�
�
�l�d�,�[Ͽ�&����P��h=�����3�8�d�u�'�.��������l��h��*���4�
�<�
�$�,�$���ǹ��^9��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����U�� G�����u�u�u�u�w�}�Wϼ��ӓ�P��S_��Hʳ�
�
�l�f�&�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�f�|�#�8�W���Y���F���*ߊ�`�l�1�u�j�4�(���H����l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�7�3�b�l�Aց�H���Z��g1����_�u�u�u�w�1��ԜY���F�N�����d�c�
�d�k�}�/���!����k>��o6��-���������L���Y�������U���u�0�1�%�8�8��Զs���K��B��*���l�"�d�4�$�:�W�������K��N�����`�d�c�
�2���������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;�b�;�(��K������D�����
��&�m�1�0�@���	����l��F1��*���
�&�
�|�w�}�������F���]���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U���}�0�<�6�9�h����L�ԓ�F�V�����
�#�
�|�~�2�W���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���M����lU�G�����_�u�u�u�w�}�W���&ƹ��_��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(ځ�L�ߓ�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���Yӄ��lS��\�����4�1�0�&�w�`����K����T9�� Y��U���u�:�;�:�g�f�}���Y����F ��h_�E���e�4�1�0�$�}����Ӗ��P��N����u� �
�
�a�m��������@��V�����'�6�o�%�8�8�ǿ�&����P��h=�����3�8�c�u�'�.��������l��1����y�4�
�<��.����&����U��B�����2�6�0�
��.�F߁�
����9F����ߊu�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���H����lW��N�����u�u�u�u�w�}����L����9��1�����&�u�h�4��2�����ғ�T�_�����:�e�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��^�����|�u�=�;�]�}�W���Y���Q��1�Gڊ�
�
�1�'�$�l�K���	����@��AX��G��x�d�1�"�#�}�^�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����`�d�g�
������
���F��h�����#�a�d�g�z�l��������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�7�3�b�l�E߁�&ù��W��D_��Hʴ�
�:�&�
�!�i�G��T����\��XN�N���u�u�u�0�$�}�W���Y���F��B��*��e�0�e�4�3�8����D�Ĕ�]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u� �
�
�a�m��������@��YN�����&�u�x�u�w�?����H����V9��T�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�l����K��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Eށ�
����O�C��U���u�u�u�u�w�?����H����V9��T�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�?����H����V9��T�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����d�g�
�
��8�W�������A	��D�X�ߊu�u� �
��k�G���I����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�b�3�8�a�}��������B9��h��D���8�d�y�4��4�(�������@��Q��M���%�&�2�6�2��#���Hù��^9��=N��U���<�_�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��m�^ϱ�Y�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��hV��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�e�3�:�d�^�������9F�N��U���u� �
�
�a�m�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u� �
�
�a�m�������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���Tӄ��lS��\�����1�u�&�<�9�-����
���9F���*ߊ�c�e�0�e�3���������PF��G�����<�
�4�2���(������]�� 1��G���;��;�0�`�8�C�������T��h��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�f�����I�ƭ�l��h�����
�!�
�&��q��������V��c1��Dڊ�&�
�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���d�3�8�d�~�}����s���F�N�����`�d�g�
���F��Y����R��hY��*��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��hW��U���;�_�u�u�w�}�W�������P��h��*��i�u�;��9�8�@���M���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�`�d�e��(߁�H���Z��V ��*݊�
�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��C���!�0�u�u�w�}�W���Yӄ��lS��\�����1�u�h�<��<����&����9F�N��U���0�_�u�u�w�}�W�������P��h��*��i�u�����/���!����k>��o6��-�����n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������lW��1��E���d�4�&�2�w�/����W���F�U��@��g�
�
�
�2���������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;�c�;�(��H������D�����
��&�d��.�(��Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�*���
�|�u�u�5�:����Y�����F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����4�
�:�&��+�(���Y����P	��1��*���d�%�|�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�l�|�~�)����Y���F�N�� ���
�c�e�0�g�*�F��Y����\��h�����n�u�u�u�w�8����Y���F�N�� ���
�c�e�0�g�*�F��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�5�;�B��Kù��9��S�����h�!�%�g��8�(��N���W��X����n�_�u�u�z�?����H����V9��V
�����u�&�<�;�'�2����Y��ƹF��B��*��e�0�d�4�3�8�ށ�
����l��TN����0�&�4�
�>�����*����9��Z1�U���&�2�6�0��	���&����V�V�����&�$��
�#�����UӇ��@��T��*���&�d�
�&��t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�d�1�0�F���Y����l�N��U���u�7�3�`�f�o�(���&����V��R�����:�&�
�#�c�n�E��Hӂ��]��G�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���I����l_����ߊu�u�u�u�w�}����&����l��h�����d�i�u�%�4�3����Oǹ��F�N�����u�|�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y�Ʈ�U9��X�*���
�1�'�&�f�a�W�������l
��1�G���d�1�"�!�w�t�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����d�g�
�
��9����H���R��X ��*���a�e�g�x�f�9� ���Y����F�N�����u�u�u�u�w�}�Wϼ��ӓ�T��R1�����0�&�u�h�u��L���Y�������U���u�0�1�%�8�8��Զs���K��B��*��e�0�d�6�g�<����Y����V��C�U���7�3�`�d�e��(ށ�ù��@��h����%�:�0�&�6�����	����l��F1��*���d�3�8�g�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��m�^������F�N��U���7�3�`�d�e��(ށ������T�����2�6�d�_�w�}�W������F�N��U���7�3�`�d�e��(ށ������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����9��^��*ۊ�0�u�&�<�9�-����
���9F���*ߊ�c�e�0�d�4�l��������\������}�%�6�y�6�����
����g9�� 1����u�%�&�2�4�8�(���
����U��^����<�
�&�$���ց�
������D�����
��&�d��.�(���Y����V��=N��U���u�3�}�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��_�����e�|�:�u��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�d����A����AF�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����l�|�|�!�2�}�W���Y���F��B��*��e�0�d�6�f�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��e�0�d�6�f�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�5�;�B��Kù��9�������%�:�0�&�w�p�W�������lW��1��D���
�&�<�;�'�2�W�������@N��h<�����
�
�y�<��<����&������e�����0�`�u�;��3�������R��^	������
�!�
�$��[Ͽ�&����P��h=����
�&�
�e�w�-��������`2��CW�����y�4�
�<��.����&����l ��hW��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�=�;�_�w�}�W���Y�Ʈ�U9��X�*���
�d�i�u�9�����N����l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�m����@����[��=N��U���u�u�u� ���A����ד�F���'���0�b�0�`�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��Q1��D��
�
�
�d�k�}��������l��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���؁�
����F��R ��U���u�u�u�u�5�;�B��Kù��9��R�����4�2�
�
��f�W���Y����_��=N��U���u�u�u� ���A����ד�F�L��-���������/���!����k>��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�h�F��&����D��V�����'�6�&�{�z�W�W�������P��h��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������F��^�����3�
�`�d�'�q��������V��c1��Dۊ�&�
�e�u�'�.��������l��h��*���4�
�<�
�$�,�$����֓�@��d��Uʷ�2�;�u�u�w�}����Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���'�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ�ӈ��N��h�����#�
�u�u�/�)����&����P��G\��\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�l�3�:�e�^ϱ�Y�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���Yӄ��lS��\�����"�d�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���Yӄ��lS��\�����"�d�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʷ�3�`�d�m��9����	����P��G]��Hʴ�
�:�&�
�!�i�G��T����\��XN�N���u�7�3�`�f�e�(�������Z�C��Aۊ� �g�d�
�f�l�Z������\F��dךU���x�7�3�`�f�e�(���������^	�����0�&�u�x�w�}����L����9��S��ۊ�&�<�;�%�8�}�W�������Q��1�Mފ�1�'�'�2�e�h�[Ͽ�&����P��h=����
�&�
�b�w�-��������`2��C\�����g�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�w�5��ԜY���F�N�����d�m�
�1�%�.�F��Y����\��h��A��d�x�d�1� �)�W���s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�m�3�:�o�^������F�N��U���7�3�`�d�o�����
���F��Q1��D��
�1�'�'�0�o�B��Y���F��[�����u�u�u�u�w�(�(ځ�A�ғ�W��D�I����n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϼ��ӓ�^��T����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��V�*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&���� W�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ԓ�@��G��U���;�_�u�u�w�}�W�������^��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}����&����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��B��*��a�6�d�4�$�:�W�������K��N�����`�d�m�
�2���������PF��G�����4�
�0�u�'�.��������l��1����y�4�
�<��.����&����l ��h\����u�0�<�_�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�e�����A�����YNךU���u�u�u�u�"��(��M����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u� �
��e�C���H���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������lW��1��U���<�;�%�:�2�.�W��Y����F ��h_�A���
�&�<�;�'�2�W�������@N��h'��0����0�8�b��8�(��L�ƭ�l��h�����
�!�m�3�:�o�[ϲ�&ƹ��^��B�����2�6�0�
��.�Eց�
����l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���Kʹ��^9��G�����_�u�u�u�w�}�W���&ƹ��R��N�U�������#�/�(�������V��=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�Eׁ�
����O��_�����u�u�u�u�w�(�(ځ�A�ғ�F���@��m�
�d�_�w�}�W������F�N��U���7�3�`�d�o��F��YѾ��k>��o6��-���������/���!��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�m�a� �l�����Ƽ�\��D@��X���u�7�3�`�f�e�(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�g�y�6�����
����g9��W�����m�_�u�u�2�4�}���Y���Z �F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��GҊ�&�
�b�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����^�G�����_�u�u�u�w�}�W���&ƹ��R��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(ځ�A�ғ�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���Yӄ��lS��]�����4�1�0�&�w�`����K����T9�� Y��U���u�:�;�:�g�f�}���Y����F ��h\�D���e�4�1�0�$�}����Ӗ��P��N����u� �
�
�n�l��������@��V�����'�6�o�%�8�8�ǿ�&����P��h=�����3�8�c�u�'�.��������l��1����y�4�
�<��.����&����U��B�����2�6�0�
��.�F߁�
����9F����ߊu�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���H����lW��N�����u�u�u�u�w�}����L����9��1�����&�u�h�4��2�����ғ�T�_�����:�e�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��^�����|�u�=�;�]�}�W���Y���Q��1�Fۊ�
�
�1�'�$�l�K���	����@��AX��G��x�d�1�"�#�}�^�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����`�g�f�
������
���F��h�����#�a�d�g�z�l��������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�7�3�b�o�Dށ�&ù��W��D_��Hʴ�
�:�&�
�!�i�G��T����\��XN�N���u�u�u�0�$�}�W���Y���F��B��*��d�0�e�4�3�8����D�Ĕ�]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u� �
�
�n�l��������@��YN�����&�u�x�u�w�?����K����V9��T�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�l����K��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Eށ�
����O�C��U���u�u�u�u�w�?����K����V9��T�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�?����K����V9��T�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����g�f�
�
��8�W�������A	��D�X�ߊu�u� �
��d�F���I����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�b�3�8�a�}��������B9��h��D���8�d�y�4��4�(�������@��Q��M���%�&�2�6�2��#���Hù��^9��=N��U���<�_�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��m�^ϱ�Y�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��hV��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�e�3�:�d�^�������9F�N��U���u� �
�
�n�l�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u� �
�
�n�l�������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���Tӄ��lS��]�����1�u�&�<�9�-����
���9F���*ߊ�l�d�0�e�3���������PF��G�����<�
�4� �;�2����&�ԓ�lV�^ �����9�:�!�:��o���Y����R��[-�����
�g�0�a�w�3�:�������G��h_����u�%�&�2�4�8�(���
�ѓ�@��N��*���
�&�$���)�F���������D�����
��&�l�1�0�O���	����l��F1��*���e�3�8�l�]�}�W������F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��m�^Ϫ���ƹF�N��U��� �
�
�l�f�8�G���Y���[��Y1������;�'�9�f��(������@[�I����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���Hù��^9��N�����u�u�u�u�w�}����L����9��1��U��}�h�<�
�6�(��������T��h^����'�h�r�r�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��L���8�m�|�!�2�}�W���Y���F��B��*��d�0�e�1�w�`�_������]��t�����d�
�
�y�8�5���^���9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�`�;���PӒ��]FǻN��U���u�u� �
��d�F���I����[�S�����;�4��;�%�1�F݁�&����G��DS�X���_�u�u�u�w�1��ԜY���F�N�����g�f�
�
��l�K���!��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�l�d�2�m� ������]F��X�����x�u�u�7�1�h�E��&����D��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�
�$��[ϻ�����WR��B1�Cۊ�g�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�f�����P�����^ ךU���u�u�3�}��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�F�������F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��B���8�c�u�;�w�2�_ǿ�&����G9��1�Hʰ�<�6�;�a�1��B���	���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�G������O��_�����u�u�u�u�w�(�(ځ�@�ד�lV��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(ځ�@�ד�lV��R_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s�����h[��L���0�d�4�1�2�.�W������ 9��P1�B���u�u�u�:�9�2�G��s���K��B��*��d�0�d�4�3�8����
������T��[���_�u�u� ���N����ד�W��D�����2�
�'�6�m�-����
ۇ��@��T��*���&�b�3�8�a�}��������B9��h��D���8�d�y�4��4�(�������@��Q��M���%�&�2�6�2��#���Hù��^9��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������lT��1��D���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Dڊ�&�
�|�u�?�3�}���Y���F�U��@��f�
�
�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�`�g�d��(ށ�����@W�
N��*���&�
�#�a�f�o�Z������\F��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���؁�
����F��R ��U���u�u�u�u�5�;�B��J¹��9��S�����h�4�
�:�$�����I���W��X����n�u�u�u�w�8����Y���F�N�� ���
�l�d�0�f�<����
���D��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u� ���N����ד�VV��D��ʥ�:�0�&�u�z�}�Wϼ��ӓ�
U��R1�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���K¹��^9��G�����u�u�u�u�w�}�Wϼ��ӓ�
U��R1����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�Wϼ��ӓ�
U��R1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʷ�3�`�g�f���(���Y����T��E�����x�_�u�u�"��(��H����l��h�����%�:�u�u�%�>����	������D�����
��&�b�1�0�A���	����l��F1��*���d�3�8�d�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1����u�0�<�_�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��C���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��PӉ��N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��h��*���u�'�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�g�;���P����[��=N��U���u�u�u� ���N����ד�VW�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u� ���N����ד�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h[��L���0�d�1�u�$�4�Ϯ�����F�=N��U���
�
�l�d�2�l�ށ�
����l��TN����0�&�<�
�6�(��������T��h_����4� �9�:�#�2�(������Z��V �����!�:�
�g�2�h�W���4����_%��C��*���0�b�u�%�$�:����&����GQ��D��Yʴ�
�<�
�&�&��(���H����lW�������6�0�
��$�d����A�ƭ�l��h�����
�!�e�3�:�d�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u� �
��d�F���H����[��Y1������;�'�9�f��(��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��t�W������F�N��Uʷ�3�`�g�f���(��E�ƥ�l+��B�����:�
�g�0�f�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:��ӊ�&�
�|�u�?�3�}���Y���F�U��@��f�
�
�
�f�a�W���4����_%��C��*���0�`�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y�Ʈ�U9��W�*���
�d�i�u�9�����:����\
��1��B�ߊu�u�u�u�;�8�}���Y���F�U��@��f�
�
�
�f�a�W͆�!����k>��o6��-���������/��Y���F��Y
�����u�u�0�1�'�2����s���F���*ߊ�l�d�0�d� �l�����Ƽ�\��D@��X���u�7�3�`�e�n�(���&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�
�&�
�{�8�����ғ�F9��_��G���%�&�2�6�2��#���H¹��^9��N��*���
�&�$���)�(���&����C9��P1������&�d�
�$��^���Yӄ��ZǻN��U���3�}�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�f�;���P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9�� 1����u�;�u�:��<�(���
����9��
N�����;�a�3�
�b�l����PӉ��N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��h��*���u�'�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�g�;���P����[��=N��U���u�u�u� ���N����ד�VW�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u� ���N����ד�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h[��Eߊ�
�
�1�'�$�m�����Ƽ�\��D@��X���u�7�3�`�d�h��������@��V�����'�6�o�%�8�8�ǿ�&����P��h=����
�&�
�d�w�-��������`2��C_�����d�y�4�
�>�����*����R��D��F���%�&�2�6�2��#���Hƹ��^9��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����9��1��E���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Dފ�&�
�f�|�#�8�W���Y���F���*ߊ�e�
�
�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�f�1�0�F���Y����l�N��U���u�7�3�`�d�h��������@��S�����;�!�9�c��u�W���Y����G	�UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����W����ߊu�u�u�u�w�}����&����V9��V
�����u�h�4�
�8�.�(���M���K�
�����e�n�u�u�w�}����Y���F�N��U���
�
�e�
������
���F��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�h�D����֓�W��D����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��^�����4�1�0�&��.����	����	F��X��¡�%�'�2�g�a�q��������V��c1��D؊�&�
�d�u�'�.��������l��h��*���!�%�g�
�"�l�Gށ�H���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�F݁�
����O��_�����u�u�u�u�w�(�(ځ�Iƹ��9��S�����h�!�%�g��(�F��&���K�
�����e�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��G���!�0�u�u�w�}�W���Yӄ��lS��[��*ڊ�1�'�&�d�k�}��������P�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�g��(߁�����@W�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����J�ӓ�lV��R^�����;�%�:�0�$�}�Z���Yӄ��lS��[��*ڊ�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���H����^9��N��*���
�&�$���)�D���������D�����
��&�d��.�(��Y����Z��D��&���!�`�3�8�f�t�W�������9F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�g�1�0�F���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�f�����J����AF�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�|�u�?�3�}���Y���F�U��@��`�0�e�6�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��&����P��V�����'�6�&�{�z�W�W������� V��R1�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������J��G1�����0�
��&�d�;���s���Q��Yd��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�u�?�3�}���Y���F�U��@��`�0�e�6�f�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��&����WW��D��ʥ�:�0�&�u�z�}�Wϼ��ӓ�S��h^��D���&�2�
�'�4�g��������Q9��^�����$�y�4�
�>�����*����T��D��D���%�&�2�6�2��#���J����lT�N�����;�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��_��U���;�_�u�u�w�}�W������� V��R1�����h�4�
�:�$�����I���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�`�f�b�8�G���Y����Q9��^�����$�n�u�u�w�}����Y���F�N��U���
�
�e�
���F��YѾ��k>��o6��-���������/���!��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�e�
������
������T��[���_�u�u� ���Gځ�&ù��9��D��*���6�o�%�:�2�.�����ƥ�l��R��*���1�'�4�
�"�o�C���UӇ��@��T��*���&�d�
�&��l�W������� 9��h_�L���y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� 9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��F����Ƣ�GN��Y1�����e�'�4�
�2�9����@ǹ��[��G1�����9�d�e�|�6�9�_�������l
��h^��U���!�:�1�
�"�l�Oց�K�����YNךU���u�u�u�u�"��(��&����D��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�7�1�h�D����֓�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h[��Eߊ�
�
�1�'�$�m�����Ƽ�\��D@��X���u�7�3�`�d�h��������@��V�����'�6�o�%�8�8�ǿ�&����P��h=����
�&�
�d�w�-��������`2��C_�����d�y�4�
�>�����*����R��D��F���%�&�2�6�2��#���Hƹ��^9��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����9��1��D���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Dފ�&�
�f�|�#�8�W���Y���F���*ߊ�e�
�
�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�f�1�0�F���Y����l�N��U���u�7�3�`�d�h��������@��S�����;�!�9�c��u�W���Y����G	�UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����W����ߊu�u�u�u�w�}����&����V9��V
�����u�h�4�
�8�.�(���M���K�
�����e�n�u�u�w�}����Y���F�N��U���
�
�e�
������
���F��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�h�D����ד�W��D����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��^�����4�1�0�&��.����	����	F��X��¡�%�'�2�g�a�q��������V��c1��D؊�&�
�d�u�'�.��������l��h��*���!�%�g�
�"�l�Gށ�H���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�F݁�
����O��_�����u�u�u�u�w�(�(ځ�Iƹ��9��S�����h�!�%�g��(�F��&���K�
�����e�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��G���!�0�u�u�w�}�W���Yӄ��lS��[��*ۊ�1�'�&�d�k�}��������P�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�g��(ށ�����@W�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����J�ӓ�lW��R^�����;�%�:�0�$�}�Z���Yӄ��lS��[��*ۊ�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���H����^9��N��*���
�&�$���)�D���������D�����
��&�d��.�(��Y����Z��D��&���!�`�3�8�f�t�W�������9F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�g�1�0�F���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�f�����J����AF�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�|�u�?�3�}���Y���F�U��@��`�0�d�6�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��&����P��V�����'�6�&�{�z�W�W������� V��R1�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������J��G1�����0�
��&�d�;���s���Q��Yd��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�u�?�3�}���Y���F�U��@��`�0�d�6�f�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��&����WW��D��ʥ�:�0�&�u�z�}�Wϼ��ӓ�S��h_��D���&�2�
�'�4�g��������Q9��^�����$�y�4�
�>�����*����T��D��D���%�&�2�6�2��#���J����lT�N�����;�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��_��U���;�_�u�u�w�}�W������� V��R1�����h�4�
�:�$�����I���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�`�f�b�8�F���Y����Q9��^�����$�n�u�u�w�}����Y���F�N��U���
�
�e�
���F��YѾ��k>��o6��-���������/���!��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�e�
������
������T��[���_�u�u� ���Gځ�&¹��9��D��*���6�o�%�:�2�.�����ƥ�l��R��*���1�'�4�
�"�o�C���UӇ��@��T��*���&�d�
�&��l�W������� 9��h_�L���y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� 9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��F����Ƣ�GN��Y1�����e�'�4�
�2�9����@ǹ��[��G1�����9�d�e�|�6�9�_�������l
��h^��U���!�:�1�
�"�l�Oց�K�����YNךU���u�u�u�u�"��(��&����D��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�7�1�h�D����ד�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h[��Eߊ�
�
�1�'�$�m�����Ƽ�\��D@��X���u�7�3�`�d�h��������@��V�����'�6�o�%�8�8�ǿ�&����P��h=����
�&�
�d�w�-��������`2��C_�����d�y�4�
�>�����*����R��D��F���%�&�2�6�2��#���Hƹ��^9��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����9��1��G���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Dފ�&�
�f�|�#�8�W���Y���F���*ߊ�e�
�
�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�f�1�0�F���Y����l�N��U���u�7�3�`�d�h��������@��S�����;�!�9�c��u�W���Y����G	�UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����W����ߊu�u�u�u�w�}����&����V9��V
�����u�h�4�
�8�.�(���M���K�
�����e�n�u�u�w�}����Y���F�N��U���
�
�e�
������
���F��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�h�D����ԓ�W��D����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��^�����4�1�0�&��.����	����	F��X��¡�%�'�2�g�a�q��������V��c1��D؊�&�
�d�u�'�.��������l��h��*���!�%�g�
�"�l�Gށ�H���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�F݁�
����O��_�����u�u�u�u�w�(�(ځ�Iƹ��9��S�����h�!�%�g��(�F��&���K�
�����e�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��G���!�0�u�u�w�}�W���Yӄ��lS��[��*؊�1�'�&�d�k�}��������P�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�g��(݁�����@W�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����J�ӓ�lT��R^�����;�%�:�0�$�}�Z���Yӄ��lS��[��*؊�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���H����^9��N��*���
�&�$���)�D���������D�����
��&�d��.�(��Y����Z��D��&���!�`�3�8�f�t�W�������9F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�g�1�0�F���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�f�����J����AF�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�|�u�?�3�}���Y���F�U��@��`�0�g�6�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��&����P��V�����'�6�&�{�z�W�W������� V��R1�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������J��G1�����0�
��&�d�;���s���Q��Yd��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�u�?�3�}���Y���F�U��@��`�0�g�6�f�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��B��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��&����WW��D��ʥ�:�0�&�u�z�}�Wϼ��ӓ�S��h\��D���&�2�
�'�4�g��������Q9��^�����$�y�4�
�>�����*����T��D��D���%�&�2�6�2��#���J����lT�N�����;�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��_��U���;�_�u�u�w�}�W������� V��R1�����h�4�
�:�$�����I���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�`�f�b�8�E���Y����Q9��^�����$�n�u�u�w�}����Y���F�N��U���
�
�e�
���F��YѾ��k>��o6��-���������/���!��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�e�
������
������T��[���_�u�u� ���Gځ�&����9��D��*���6�o�%�:�2�.�����ƥ�l��R��*���1�'�4�
�"�o�C���UӇ��@��T��*���&�d�
�&��l�W������� 9��h_�L���y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� 9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��F����Ƣ�GN��Y1�����e�'�4�
�2�9����@ǹ��[��G1�����9�d�e�|�6�9�_�������l
��h^��U���!�:�1�
�"�l�Oց�K�����YNךU���u�u�u�u�"��(��&����D��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�7�1�h�D����ԓ�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���Yӄ��lS��^��*ڊ�1�'�&�e�k�}����J����lT�� F�X��1�"�!�u�~�W�W���T�Ʈ�U9��_�����4�1�0�&�w�.����	����@�CךU��� �
�
�d���(�������l��^	�����u�u�'�6�$�u��������B9��h��*���
�y�4�
�>�����*����W��D��E���%�&�2�6�2��#���@����l^�V�����&�$��
�#�m����@���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�Fށ�
����O��_�����u�u�u�u�w�(�(ځ�Hù��9��S�����h�4�
�:�$�����J���W��X����n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����V��D��\���=�;�_�u�w�}�W���Y����9��1��E���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��L���8�m�|�!�2�}�W���Y���F��B��*��
�
�
�1�%�.�F��Y����\��h��A��g�x�d�1� �)�W���s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��Uʷ�3�`�l�e�2�m��������[��G1�����9�c�
�}�w�}�W������]ǻN��U���9�0�_�u�w�}�W���Y����9��1��E���1�0�&�u�j��/��Y���F��Y
�����u�u�0�1�'�2����s���F���*ߊ�d�
�
�
�2�}����Ӗ��P��N����u� �
�
�f��(߁�ù��@��h����%�:�0�&�6�����	����l��F1��*���g�3�8�g�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^������F�N��U���7�3�`�l�g�8�G���I���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U��� �
�
�d���(���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z�������
W��R1����4�&�2�u�%�>���T���F��Q1��L���0�e�6�d�6�.���������T��]���6�y�4�
�>�����*����9��Z1�U���&�2�6�0��	���&����V�V�����&�$��
�#�����UӇ��@��T��*���&�d�
�&��t�W�������9F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����W��D��E���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�l�1�0�O������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��L���|�!�0�u�w�}�W���Y����F ��hW�*���
�0�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ʈ�U9��_�����6�d�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�7�3�`�n�m�����ƭ�@�������{�x�_�u�w�(�(ځ�Hù��9��h�����%�:�u�u�%�>��������]��h��Yʼ�
�4�;�
���[Ϸ�&����@9��R1�U����<�&�a�2�k�W���
����@��d:��݊�&�
�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
�ߓ�@��N��*���
�&�$���)�G������F�U�����u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����V����ߊu�u�u�u�w�}����&����V9��S_��Hʼ�
�4�;�
���L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�~�}����s���F�N�����`�l�e�0�g�9�W������Z��1��A�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ߓ�@��G�����_�u�u�u�w�}�W���&ƹ��9��1��U��<�
�4�;���(��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�b�3�8�a�t����Y���F�N��U���
�
�d�
���F��Y����R��hZ��*��u�u�u�u�2�.�W���Y���F���*ߊ�d�
�
�
�f�a�W͆�!����k>��o6��-���������/��Y���F��Y
�����u�u�0�1�'�2����s���F���*ߊ�d�
�
�
�2�}����Ӗ��P��N����u� �
�
�f��(߁�¹��@��h����%�:�0�&�6�����	����l��F1��*���
�&�
�y�2�4����M����S��h�U���&�2�6�0��	���&����V�V�����&�$��
�#�����UӇ��@��T��*���&�d�
�&��t�W�������9F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�d�1�0�F���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��C���;�u�:�}�6�����&����F�R�����a�3�
�`�f�-�^������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����G_��D��\���'�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�e�1�0�N���PӒ��]FǻN��U���u�u� �
��l�(���&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�7�3�`�n�m�������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�Wϼ��ӓ�V��h_�����&�e�i�u�:��D�������N��N����!�u�|�_�w�}�Z�������
W��R1�����0�&�u�&�>�3�������KǻN�� ���
�d�
�
��9����H����Z��G��U���'�6�&�}�'�.��������l��h��*���4�
�<�
�$�,�$����ד�@��B�����2�6�0�
��.�N������R��^	������
�!�e�1�0�N�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����I����[��=N��U���u�u�u� ���F߁�&¹��W��D_��Hʴ�
�:�&�
�!�i�D��T����\��XN�N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����֓�@��G�����_�u�u�u�w�}�W���&ƹ��9��1�����&�u�h�4��2�����ғ�T�_�����:�e�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y����F ��hW�*���
�1�'�&�f�a�W�������l
��1�G���d�1�"�!�w�t�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����l�e�0�d�6�9����Y����C9��Y����
�}�u�u�w�2����I��ƹF�N�����_�u�u�u�w�}�W���&ƹ��9��1�����&�u�h�w��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h[��Dڊ�
�
�0�u�$�4�Ϯ�����F�=N��U���
�
�d�
���߁�
����l��TN����0�&�4�
�2�}��������B9��h��G���8�g�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�}����s���F�N�����`�l�e�0�f�>�G��Y����\��h�����n�u�u�u�w�8����Y���F�N�� ���
�d�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}����&����V9��T����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��_�����6�d�4�&�0�����CӖ��P�������4�
�<�
�$�,�$���Ĺ��^9�������6�0�
��$�l�(���&���R��^	������
�!�
�$��[Ͽ�&����P��h=����
�&�
�|�w�}�������F���]���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ד�@��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�l�3�8�o�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��G��\ʡ�0�u�u�u�w�}�W�������l_��h��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W�������
W��R1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʷ�3�`�l�e�2�l����
������T��[���_�u�u� ���F߁�&¹��l��^	�����u�u�'�6�$�u��������l��N��*���;�
�
�
�{�4�(�������V9����2���&�a�0�b�w�-��������`2��CY�����y�4�
�<��.����&����l ��h_�U���&�2�6�0��	��������F��h��*���$��
�!�g�;���s���Q��Yd��U���u�<�u�}�'�>��������lW������6�0�
��$�l�(���&�����YNךU���u�u�u�u�"��(��&����WW�
N��*���;�
�
�
�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Dڊ�&�
�|�u�?�3�}���Y���F�U��@��e�0�d�1�w�`��������9��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�(�(ځ�Hù��9��R�����4�;�
�
��f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�c�|�#�8�W���Y���F���*ߊ�d�
�
�
�f�a�W���>����lR��h_�U���u�u�0�&�w�}�W���Y�����h[��Dڊ�
�
�d�i�w��/���!����k>��o6��-��������f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h[��Dڊ�
�
�0�u�$�4�Ϯ�����F�=N��U���
�
�d�
���ށ�
����l��TN����0�&�4�
�2�}��������B9��h��*���
�y�0�<�4�3�C���&����l�������6�0�
��$�l�(���&���R��^	������
�!�
�$��[Ͽ�&����P��h=����
�&�
�|�w�}�������F���]���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�f�t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����:�}�4�
�8�.�(���&���V��T��A���
�`�d�%�~�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ߓ�@��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�t�^Ϫ���ƹF�N��U��� �
�
�d���(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʷ�3�`�l�e�2�l� ��E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�?����@�ߓ�W��P�����a�
�f�i�w�-��������9��N�Dʱ�"�!�u�|�]�}�W���&ƹ��
9��S�����h�!�%�g��(�F��&���K�
�����e�n�_�u�w�p����L����l��E��Dʴ�&�2�u�'�4�.�Y��s���Q��1�L���1�0�&�
�$�4��������C��R�����`�l�l�4�3�����M���R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�`�u�'�.��������l��h��*���4�
�<�
�$�,�$���ƹ��^9��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�Wϼ��ӓ�_��S
����i�u�%�6�9�)���&����F��S�����|�_�u�u�w�}����Y�έ�l��D�����
�u�u�%�$�:����&����GS��D��\���=�;�_�u�w�}�W���Y����9��1�����&�u�h�4��2�����ғ�T�_�����:�e�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y����F ��hW�*���'�&�d�i�w�-��������9��N�Dʱ�"�!�u�|�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��Q1��L���4�1�0�&�w�`����L����l��E1����f�n�u�u�w�}����Y���F�N��U���
�
�`�
�3�/���E����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�7�3�`�n�d�������]F��X�����x�u�u�7�1�h�N����֓�@��Y1�����u�'�6�&��-�������T9��R��!���d�
�&�
�a�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�b�3�:�l�^�������9F�N��U���u� �
�
�b�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����`�l�l�6�g�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�5�;�B��@������^	�����0�&�u�x�w�}����L����l��h�����%�:�u�u�%�>����	������D�����
��&�g�1�0�F���	����l��F1��*���
�&�
�y�6�����
����g9��1����u�%�&�2�4�8�(���
�ӓ�@��d��Uʷ�2�;�u�u�w�}����Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h_��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�`�3�8�c�t�^Ϫ���ƹF�N��U��� �
�
�`��8�W������]��[����_�u�u�u�w�1��ԜY���F�N�����l�l�6�d�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�h�N����ƭ�@�������{�x�_�u�w�(�(ځ�Lʹ��l��^	�����u�u�'�6�$�u����&����J��Y1��*؊�
�y�<�
��o���Y����e9��R1�U���&�2�6�0��	��������F��h��*���$��
�!��.�(������T9��R��!���a�3�8�f�w�-��������`2��C[�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��Q1��L���1�u�h�<���E���J���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�`�l�n�9�W������lT��h\�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&���� O�C��U���u�u�u�u�w�?����@�ߓ�F���%���
�
�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y����F ��hW�*��i�u�;����(��Y���F��[�����u�u�u�u�w�(�(ځ�Lʹ��Z�6��-���������/���!����k>��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u� ���Bց��ƭ�@�������{�x�_�u�w�(�(ځ�Lʹ��9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��q��������l ��[�*��u�%�&�2�4�8�(���
�Г�@��N��*���
�&�$���)�(���&����C9��P1������&�`�3�:�i�}���Y����]l�N��Uʼ�u�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�c�1�0�B������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��D��\ʴ�1�;�!�}�/�)����&����R��G\��U���6�;�!�9�f�m�^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�`�3�:�i�^�������9F�N��U���u� �
�
�b�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����`�l�l�"�f�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�6�
���2�������V9��Q��D���%�u�h�_�w�}�W�������u	��{��*���0�d�'�2�e�m�W����ο�_9��G]�����2�g�a�}�~�`�P���Y����l�N��Uʦ�9�!�%�l�>�;�(��@����9F������1�
� �g�o��E��Y���D��F��*���
�a�f�h�6�����&����O��[��W���_�u�u�-�#�2�݁�����9��R��W���"�0�u�<��4�1���5����@9��P1�B���u�%�6�;�#�1�D��Y����D��d��Uʰ�<�6�;�f�1��B���	���D�������d�'�2�d�a�}�W�������l
��hZ�����u�e�n�u�w�8�����ғ�F9��_��G��u�d�u�=�9�u��������V��_�����2�d�a�u�w�-��������lT�R��U��n�u�u�0�>�>��������T��N�U��u�=�;�}��8�(��A����C9��Y�����a�u�9�0�u��}���Y����P	��h��G��
�g�i�u�f�}����Q�Փ�V��W�Hʴ�
�:�&�
�!��^ϻ�
���]ǻN��&������!�f�k����H�ד� F�d��U���u�4�
�:�$�����Iӑ��]F��Z��B���2�g�c�}�~�`�P���Y����l�N��Uʲ�%�3�
�`�b�-�L���YӀ��`#��t:�����
� �d�g��n�K���Y���F��B��*��d�0�d�$�w�5��������_��h��*��e�u�u�d�~�8����Y���F��B��*��f�0�g�$�l�}�Wϸ�&����}"��C��*���3�
�l�d�'�}�Jϼ��ӓ�V��h_��E�ߊu�u��!�%�l�F���H����W��h�I���u�u�u�u�4���������C9��h��*���
�c�m�"�2�}����MŹ��lT��1��]���h�r�r�u�;�8�}���Y���U5��r"��!���
�c�'�2�e�l�L���YӀ��G��1�G���3�
�d�e�'�}�J�ԜY���F��h��3����:�
�l�2�l����K����D��F����
�0�
�b�d�m�W���H����_��=N��U���u��������&����Q��d��Uʳ�
���g��)�Oہ�&����^��G]��H�ߊu�u�u�u��%�"�������R��B1�Cۊ�d�"�0�u�$�1����&����lT�� 1��]���h�r�r�u�;�8�}���Y���Q��1�E���d�$�n�u�w�;�(���5�Ԣ�F��1��*��d�%�u�h�'�����&�ד�F9��W��@�ߊu�u��-��	����&�ғ�]9��G1��D���
�l�l�%�w�`��������l��C�����0�}�%�6�9�)���&����uO������%��&�9�����A¹��O��N�������g��#�e�(�������V9��h_�F���u�h�_�u�w�}�W���&����Z9��T��*���!�3�
�l�b�-�W����ο�_9��G\��*���d�c�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�
��(�F��&����F�Q��*��f�4�1�0�$�}�JϪ�	����F9�� ]��D��x�d�1�"�#�}�^�ԜY�ƪ�lS��[�����0�&�u�h�#�-�Cށ����� R�C��U���;�:�e�n�]�}�W������_��h��U���<�;�%�:�2�.�W��Y����Q9��W�*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O����ߊu�u�u�u�w�}����H����P��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�3���N������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӀ��9��]�����&�<�;�%�8�8����T��� ��1�@ي�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���J����^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h]�\���=�;�_�u�w�}�W���Y����lW��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����Q9��W�*��i�u� �
��e�C���B���F���@��`�
�0�u�$�4�Ϯ�����F�=N��U���`�d�`�
�2���������PF��G�����4�
�0�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF�F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��F���8�f�|�|�w�5��ԜY���F�N��*ߊ�l�f�"�d�k�}��������\��h_�U���u�u�0�&�w�}�W���Y��� ��1�@ي�0�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=N��U���`�f�`�0�g�<����
�����h��D���
�d�g�x�f�9� ���Y����F�Q��*��
�
�
�1�%�.�F��Y����V��R	��L��g�x�d�1� �)�W���s���K�Q��*��
�
�
�0�w�.����	����@�CךU���7�`�f�`�2�m��������]9��X��U���6�&�}�%�4�q��������V��c1��G���8�d�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�|�#�8�W���Y���F���@��`�0�e�6�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��U1��F���0�e�6�e�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�3���Gځ�&ù��F��D��U���6�&�{�x�]�}�W���L����l��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�n�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O����ߊu�u�u�u�w�}����J�ӓ�lV��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�?�B��L����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����Q9��^�����1�u�h�9���A����֓�]ǑN��X���7�`�f�`�2�m� ������]F��X�����x�u�u�3���Gځ�&ù��9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�d�3�:�n�^���Yӄ��ZǻN��U���3�}�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�f�;���P���G��d��U���u�u�u�3���Gځ�&ù��F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�3�
��m�(���&����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W����ӓ�S��h_�����&�e�i�u�:����Lǹ��T�_�����:�e�n�u�w�;�(ځ�Iƹ��9��S�����h�!�%�a��8�(��M���W��X����n�_�u�u�z�;�(ځ�Iƹ��9��N�����u�'�6�&�y�p�}���Y����lU��h��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O����ߊu�u�u�u�w�}����J�ӓ�lW��R^��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�?�B��L����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��U1��F���0�d�6�d�6�.��������@H�d��Uʳ�
�
�e�
���ށ�
����l��TN����0�&�4�
�2�}��������B9��h��D���8�f�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�e�~�}����s���F�N�����
�e�
�
��8�W������]��[����_�u�u�u�w�1��ԜY���F�N��*ߊ�e�
�
�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�7�b�n�B���H����[��C1��@��
�
�
�e�]�}�W��Y����lU��h��*���u�&�<�;�'�2����Y��ƹF��U1��F���0�d�"�d�6�.���������T��]���6�y�4�
�>�����*���� W��D��E�ߊu�u�0�<�]�}�W���Y���N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��_�����e�|�|�!�2�}�W���Y���F��U1��F���0�d�"�d�k�}��������\��h_�U���u�u�0�&�w�}�W���Y��� ��1�@���d�"�d�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���3�
�
�e���(�������Z�C�����`�a�%�}�w�}�W������]ǻN�����f�`�0�g�6�9����Y����^��1����e�}�u�u�w�2����I��ƓF�C�����f�`�0�g�4�m�����Ƽ�\��D@��X���u�3�
�
�g��(݁�ù��@��h����%�:�0�&�6�����	����l��F1��*���
�&�
�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�~�}����s���F�N�����
�e�
�
��8�W������]��[����_�u�u�u�w�1��ԜY���F�N��*ߊ�e�
�
�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�?�B��L����l�������%�:�0�&�w�p�W������� V��R1�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���J¹��^9��G�����u�u�u�u�w�}�Wϸ�&ƹ��9��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����V9��T�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��h[��Eߊ�
�
�d�i�w�)�B��@ƹ��9��dךU���x�3�
�
�g��(݁��ƭ�@�������{�x�_�u�w�?�B��L����l��h�����%�:�u�u�%�>����	������D�����
��&�f��.�(��s���Q��Yd��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�n�(���&���O��_�����u�u�u�u�w�?�B��L����l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�5�h�D����ԓ�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h��D��
�0�4�&�0�}����
���l�N�����
�`�`�6��.����	����	F��X��´�
�0�u�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����֓�@��B�����2�6�0�
��.�Eށ�
����F��h��*���$��
�!�e�;���UӇ��@��T��*���&�g�
�&��o�W���
����@��d:�����3�8�g�y�6�����
����g9��[�����a�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���N����lT�������6�0�
��$�l�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�u��������\��h_��U���&�2�6�0��	���&����Q�X�����:�&�
�:�>��W���	����l��F1��*���e�3�8�d�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ד�@��G�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�W���Q����\��h�����u�u�%�&�0�>����-���� 9��Z1�\ʺ�u�4�
�:�$�����&���R��^	������
�!�a�1�0�E�������C9��Y�����6�d�h�4��4�(�������@��h��*��u�'�}�%�4�3��������[��G1�����0�
��&�e�����L�ƣ�N��h�����:�<�
�u�w�-��������`2��C\�����g�|�:�u�6�����&����P9��
N��*���
�&�$���)�N�������O�C��U���u�u�u�u�w�:����&����l��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�2�'�;�(��L����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƫ�C9��h_�@���6�1�u�&�>�3�������KǻN����� �d�e�
�'�2����
����C��T�����&�}�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���H����lT����*���'�2�g�g�{�.����	�ד�l��h\�L���0�
�8�g������N���@��C��L���'�2�g�a�{�.����	�ѓ�l��h\�B���8�
�b�'�0�o�A������T9��R��!���g�
�&�
�d�}��������B9��h��@���8�g�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�`�}��������]��[��E��&�9�!�%�f�4����K������F��*���&�
�#�
�w�}��������Z9��P1�F���4�1�}�%�4�3����H�����h��Gӊ�
�0�
�b�f�}��������]��[��E��&�9�!�%�`�4����K������F��*���&�
�#�
�w�}����A����lT��G�����4�
�:�&��2����Y�ƭ�l��h�����
�!�a�3�:�o�^Ͽ��έ�l��D��ۊ�u�u�8�
�`�/���O���F��R ��U���u�u�u�u�0�-����L�ӓ�C��RN�U���6�;�!�9�e�l�}���Y���V
��QN��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�g�}����	����@��X	��*���u�%�&�2�4�8�(���
����U��Z��\ʡ�0�u�u�u�w�}�W�������F9��[�����0�i�u�%�4�3����K����F�N�����u�u�u�u�w�}�WϹ�	����S��h�����i�u��w�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƫ�C9��h_�@���u�&�<�;�'�2����Y��ƹF��E�� ��e�
�e�4�$�:�(�������A	��D�� ���
�`�
�e�w�-��������`2��C_�����d�y�3�
���8���LĹ��T9��X����<�
�&�$����������J��[1��*���
�:�%�g���(���&����F��h��*���$��
�!�c�;���UӀ��K+��c�����9�<�9�
�e�/���A����C9��P1������&�g�
�$��C�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����M����[��=N��U���u�u�u�'��(�F��&���F��h��9��� �
� �!�'�$�@݁�����S��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�C�������F��R ��U���u�u�u�u�0�-����L�ӓ�F������:�
�:�%�e��(݁�����U��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�F�������F��R ��U���u�u�u�u�0�-����L�ӓ�F������,� �
�b�%�:�E��B���F������}�%�6�;�#�1����H����C9��P1������&�d�
�$��@�������9F�N��U���u�'�
� �f�m�(��E�Ʈ�U9��[����u�u�u�u�2�.�W���Y���F�	��*���d�e�
�e�k�}�/���!����k>��o6��-���������L���Y�������U���u�0�1�%�8�8��Զs���K��E�� ��e�
�d�4�$�:�W�������K��N�����3�
�`�`�'���������PF��G�����4�
�<�
�$�,�$����ޓ�@�� B�� ���
�`�l�$�{�?����H����V9��F^����<�
�&�$����������J��d1��*���'�2�g�`�{�<�(���&����l5��D�*���
�f�u� ���D����֓�J��G1�����0�
��&�e�����M���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�Eځ�
����O��_�����u�u�u�u�w�/�(���H����CW�
N�����d�f�
�
��m�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���a�3�8�g�~�}����s���F�N�����3�
�`�`�'�}�Jϸ�&����9��P1�@��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h\�\ʡ�0�u�u�u�w�}�W�������F9��[��D��u� �
�
�d�n������ƹF�N�����u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u�'�
�"�l�Gځ�H���Q��1�Cӊ�e�_�u�u�w�}����s���F�N�����3�
�`�`�'�}�J���!����k>��o6��-���������/���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����
�`�a�%�w�.����	����@�CךU���'�
� �d�f��G���
����C��T�����&�}��-��$����N����lT��B�����2�6�0�
��.�E܁�
����F��h��9����!�m�
��8�(��M�ƭ�l��h�����
�!�a�3�:�o�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��h��*���$��
�!�c�;���P�Ƹ�V�N��U���u�u�2�%�1��B���	��� ��O#��!ػ� �
�a�d�%�:�E��B���F������}�%�6�;�#�1����H����C9��P1������&�g�
�$��E�������9F�N��U���u�'�
� �f�l�(��E�ƪ�l��u�����
�0�
�c�a�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��B���	���D��o6��-���������/���!����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�2�%�3��h�C���Y����T��E�����x�_�u�u�%����Hǹ��l��^	�����u�u�'�6�$�u�$���=����G9��h��*��f�u�%�&�0�>����-���� 9��Z1�Yʴ�
�<�
�&�&��(���M����lT����*ߊ�d�
�
�
�g�W�W�������F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��D�������9F�N��U���u�'�
� �f�l�(��E�ƪ�l��s����
�0�
�b�d�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�w�5��ԜY���F�N�����
�`�a�%�w�`����L����l��h����u�u�u�9�2�W�W���Y���F��G1��*���a�%�u�h�u��/���!����k>��o6��-�������u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���T��Q��@���:�6�1�u�$�4�Ϯ�����F�=N��U���
� �d�d��-��������]9��X��U���6�&�}�%�$�:����&����GT��Q��G���!�%�a�
�2��@��Y����G��1�����g�g�y�&�;�)��������lT��B�����8�g�
�
�2��@��Y����G�� 1�����g�a�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}��������B9��h��F���8�g�|�4�3�u��������EW��S�����8�g�
�
�2��@��Y������T�����d�e�h�&�;�)��������lT�� G�����:�}�4�
�8�.�(���&���@��C��E���'�2�g�f�~�t�W������F�N��Uʲ�%�3�
�`�n�2����Y����C9��Y�����a�_�u�u�w�}����Y����C9��Y�����6�d�h�4��4�(�������@��h��*��u�;�u�4��2����¹��F��[1�����<�'�2�g�e�t����Q����\��h��*���u�0�
�8�e��(���&����F��SN�����;�!�9�d�g�`��������l��R	��B��u�;�u�4��2����¹��F��[1�����<�'�2�g�c�t����Q����\��h��*���u�8�
�m�%�:�E��P����[��=N��U���u�u�u�'��(�F��&����W�
N��*���&�
�#�
�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��G؊�&�
�d�|�#�8�W���Y���F�	��*���d�d�
�%�8�8�K���	����@��A[��N���u�u�u�0�$�}�W���Y���F��E�� ��d�
�%�:�2�a�W͆�!���9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���'�
� �d�f��GϿ�
����C��R��U���u�u�2�%�1��B���	ù��@��h����%�:�0�&�6�����
����g9��\�����d�u� �
��k�G���H���� ��d+��6���!�`�
�0��j�F�������l��h\�F���0�
�8�d������N���@��C��E���'�2�g�f�{�.����	�ߓ�l��h\�D���0�
�8�f������N���R��^	������
�!�f�1�0�E������l_��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}��������B9��h��F���8�g�|�4�3�u��������EW��S�����8�g�
�
�2��@��Y������T�����d�e�h�&�;�)��������lT�� G�����:�}�4�
�8�.�(���&���@��C��E���'�2�g�f�~�t�W������F�N��Uʲ�%�3�
�`�n�-�W������#��x��@܊�0�
�b�d�]�}�W���Y����UF������!�9�2�6�f�`��������V��c1��Gي�&�
�g�u�9�}��������_��N�����!�%�d�<�%�:�E��PӇ��N��h�����#�
�u�u�2����&����T9��[�����}�%�6�;�#�1�F��Dӕ��l��W��*���
�b�d�u�9�}��������_��N�����!�%�b�<�%�:�E��PӇ��N��h�����#�
�u�u�:��O������� O����ߊu�u�u�u�w�}��������
9��R�����`�l�e�0�f�,�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�f�t����Y���F�N��U���
� �d�d��m�K�������P��h��*��_�u�u�u�w�1��ԜY���F�N�����
�`�l�%�w�`�U���!����k>��o6��-���������U�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�P�����`�l�%�u�$�4�Ϯ�����F�=N��U���
� �d�d��l��������\������}�%�&�2�4�8�(���
����U��_����`�d�g�
���G�������u	��{��*���0�e�'�2�e�d�[Ϫ�	����A��Y�Yʦ�9�!�%�d�>�/���K����V
��Z�*���0�
�b�`�w�8�(���Kʹ��A��Y�Yʦ�9�!�%�b�>�/���M����C9��P1������&�g�
�$��E�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����&�$��
�#�n����K����]�V�����
�#�
�u�w�8�(���Kʹ��A��Y�\ʴ�1�}�%�6�9�)����I����V
��Z�*���0�
�b�b�w�3�W���Qۇ��P	��C1��D��h�&�9�!�'�m��������O�N�����u�u�u�u�w�}��������_��N�U���9�
�:�
�8�-�Eց�&ù��T9��V�U���u�u�0�&�1�u�_�������l
��^��U���%�&�2�6�2��#���K����^9��N�����%�6�;�!�;�l�G��
����^��h�����b�l�u�;�w�<�(���
����9��
N�����%�e�<�'�0�o�D������R��X ��*���
�u�u�0��0�Eց�&����Q��N�����%�6�;�!�;�l�G��
����^��h�����b�b�u�;�w�<�(���
����9��
N����
�0�
�b�d�t�W������F�N��Uʲ�%�3�
�`�n�-�W������]��[�*��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h\�\ʡ�0�u�u�u�w�}�W�������F9��W��D��u� �
�
�a�m������ƹF�N�����_�u�u�u�w�}�W���&����W��G_��H���������/���!����k>��o6��-���_�u�u�u�w�3�W���Y����������n�_�u�u��1�(���&����lW��Q��C���%�u�h�&�3�1��������AN��D������9�
�:��2��������Q��E�����;�1�4�
�8�.�(���&���9F���*���d�a�
�g�k�}��������E��X�����;�1�<�'�0�l�D���Rӓ��Z��SF��*���&�
�#�
�~�f�W����ԓ�F9��[��G��u�!�
�:�>�����ۓ��Z��SF��*���
�a�d�u�w�3����ۇ��P	��C1��F��|�_�u�u�����@ǹ��Z�D�����6�#�6�:��3����ۏ��A��Z�\��� �&�2�0��-��������lW�d��Uʼ�a�3�
�g�d�-�W��
����\��h����� �&�2�0��n����H����M��Y�����4�
�:�&��+�(���B�����E�����'�4�
�0�3�;�(��&���F�
P��*���0�
�y�:�?�/�J���^��ƹF��X��*ۊ� �d�d�
�f�a�W���,����w*��R��G؊� �d�e�
�f�o�W���Y����G	�UךU���:�
�
�
�"�l�Cށ�M���C9��[\��*���d�f�
�d�d�}��������l�N�����f�3�
�c�f�-�W��	����9��Q��C���%�}�f�x�f�9� ���Y����F�[��#���3�
�c�b�'�}�JϮ�/����9��h_�F���}�e�1�"�#�}�D��Y����\��h[�� ��m�
�d�i�w�����A����P��h�G���u�u�:�;�8�m�L���Yӊ��l0��h��D��
�a�i�u��<�E�������_��F�U���;�:�g�|�]�}�W���&����U�� \�����h�%��9�����Iʹ��T��N����!�u�|�_�w�}����&����
V��GZ��Hʳ�
�� ���8���&����
V��G_��Eʱ�"�!�u�f�l�}�Wϲ�&ƹ��^��S
�����3�
�c�
�d�a�W�������l
��1�G���d�1�"�!�w�t�}���Y���_��h_�M���1�0�&�u�$�4�Ϯ�����F�=N��U���`�d�m�
�3�/��������]9��X��U���6�&�}�!�b�l�Oׁ�����V��Z�U���&�2�6�0��	���&����P�V�����&�$��
�#�e����K��ƹF��R	�����u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�1�(ځ�O�ޓ�W��D�I���%�6�;�!�;�k�(���Y����W	��C��\�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��X��U���;�_�u�u�w�}�W����ӓ�^��V
�����u�h�9�
��k�O�������T9��V�U���u�u�0�&�w�}�W���Y���
��1�MҊ�1�'�&�e�k�}�/���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*ߊ�c�m�4�1�2�.�W�������A	��D�X�ߊu�u�!�`�f�e�(�������l��^	�����u�u�'�6�$�u��������B9��h��B���8�d�y�!�'�o�(���&����F��h��*���$��
�!�o�;���UӇ��@��T��*���&�g�
�&��k�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�g��.�(��PӒ��]FǻN��U���u�u�!�`�f�e�(�������Z�C��Gي�0�
�`�b�e�p�FϺ�����O��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�O�������F��R ��U���u�u�u�u�;��(��A����A��N�U���6�;�!�9�a��_���Y�ƨ�D��^����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���HĹ��^9��G�����_�u�u�u�w�}�W���L����9��S�����h�4�
�:�$�����H���W��X����n�u�u�u�w�8����Y���F�N�����d�m�
�1�%�.�F��YѾ��l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���9�
�
�c�o�>�GϿ�
����C��R��U���u�u�9�
��k�O���I����Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�c�w�-��������`2��C\�����g�|�u�u�5�:����Y�����F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���A����lT��G�����u�u�u�u�w�}�Wϲ�&ƹ��^��R^��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�)�B��A˹��F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���_��h_�M���d�4�&�2�w�/����W���F�[��*��m�6�d�4�$�:�(�������A	��D�����y�4�
�<��.����&����l ��h_�U���&�2�6�0��	���&����Q�V�����&�$��
�#�j����K��ƹF��R	�����u�u�u�3��u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�b�~�2�W���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���KĹ��^9��G��U���;�_�u�u�w�}�W����ӓ�^��T�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�1�(ځ�O�ޓ�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���Yӊ��9��V��D��u�9����)����A����l��h\�A�ߠu�u�x�u�#�h�F��&����R��P �����&�{�x�_�w�}����H����D��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�b�1�0�E���Y����V��=N��U���u�3�}�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�j����K���F��R ��U���u�u�u�u�;��(��A����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�!�`�f�e�(���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z����ӓ�R��R1�����0�&�u�&�>�3�������KǻN�����d�a�
�
��9����I����Z��G��U���'�6�&�}�'�.��������l�� 1����y�4�
�<��.����&����l ��h\����u�0�<�_�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y����G9��V�*���
�1�'�&�g�a�W�������l
��1�G���d�1�"�!�w�t�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���b�3�8�d�~�}����s���F�N�����
�m�c�0�g�<����
�����T�����c�
�}�u�w�}�������9F�N��U���0�_�u�u�w�}�W����ӓ�R��R1�����0�&�u�h�u��L���Y�������U���u�0�1�%�8�8��Զs���K��C1��D��
�
�
�1�%�.�FϿ�
����C��R��U���u�u�9�
��e�A���I����A��1�����
�'�6�o�'�2��������T9��R��!���d�
�&�
�a�}����J����lT�� B�����2�6�0�
��.�Eׁ�
����F��h��*���$��
�!�`�;���P�����^ ךU���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�@�������F��R ��U���u�u�u�u�;��(��O����l��E��D��u�8�
�f�%�:�E��Q���F��@ ��U���_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����lW��1��E���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��D݊�&�
�c�|�#�8�W���Y���F���@��a�
�
�
�3�/���E�ƭ�l��D�����d�g�x�d�3�*����P���F�N�����u�u�u�u�w�}����&����l��h�����d�i�u��u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���_��h_�C���e�6�e�4�$�:�W�������K��N�����
�m�c�0�g�>�G���
����C��T�����&�}�%�6�{�<�(���&����l5��D�*���
�c�u�%�$�:����&����GT��Q��G���u�u�7�2�9�}�W���Yӏ��N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�O�������O�C��U���u�u�u�u�w�1�(ځ�A�Г�lV��R^��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�)�B��MŹ��9��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�[��*��c�0�e�6�f�<����Y����V��C�U���9�
�
�m�a�8�G���H����Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�c�w�-��������`2��C\�����g�y�4�
�>�����*����Q��D��C�ߊu�u�0�<�]�}�W���Y���N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��Y�����c�|�:�u��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��B���8�g�|�|�w�5��ԜY���F�N��*ߊ�m�c�0�e�4�l�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���@��a�
�
�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�!�b�l�Cف�&ù��Z�Q=����
�0�
�b�o�W�W���T�Ơ�lS��Z�����"�d�4�&�0�}����
���l�N��*ߊ�m�c�0�e� �l��������\������}�%�6�y�6�����
����g9��Y�����c�_�u�u�2�4�}���Y���Z �F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��G݊�&�
�c�|�~�)����Y���F�N�����d�a�
�
��8�W������]��[����_�u�u�u�w�1��ԜY���F�N��*ߊ�m�c�0�e� �l�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�1�(ځ�A�Г�lW��S
����4�&�2�u�%�>���T���F��h[��M���0�d�4�1�2�.�(�������A	��N�����&�4�
�<��.����&����l ��h_�U���&�2�6�0��	���&����Q�N�����;�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��Y��U���;�_�u�u�w�}�W����ӓ�R��R1�����0�&�u�h�6�����&����lT�C��U���;�:�e�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�c�|�!�2�}�W���Y���F��C1��D��
�
�
�1�%�.�G��Y����\��h��A��g�x�d�1� �)�W���s���F�R��U���u�u�u�u�w�1�(ځ�A�Г�lW��S
����i�u��w�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ơ�lS��Z�����4�1�0�&�w�.����	����@�CךU���!�`�d�a���(�������l��^	�����u�u�'�6�$�u��������B9��h��B���8�d�y�!�'�o�(���&����F��h��*���$��
�!�o�;���UӇ��@��T��*���&�g�
�&��k�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�g��.�(��PӒ��]FǻN��U���u�u�!�`�f�i�(���&����V��R�����g�
�0�
�b�j�E��Hӂ��]��G�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���A����lT��N�����u�u�u�u�w�}����&����l��h�����d�i�u�%�4�3����Oǹ��F�N�����u�|�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l�� 1����|�u�=�;�]�}�W���Y���_��h_�C���d�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����RNךU���u�u�u�u�#�h�F��&����R��R��U��w��n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������^��h��*���u�&�<�;�'�2����Y��ƹF��C1��D��
�
�
�0��.����	����	F��X��´�
�0�u�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����ޓ�@�� GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����Q��D��C���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�g��.�(��P����[��=N��U���u�u�u�!�b�l�Cف�&¹��F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�9�
��e�A���H����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����G9��V�*���
�0�u�&�>�3�������KǻN�����d�a�
�
��8�(�������A	��N�����&�4�
�0�w�-��������`2��C_�����d�y�4�
�>�����*����^��D��B���%�&�2�6�2��#���KĹ��^9��d��Uʷ�2�;�u�u�w�}����Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���'�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�m�1�0�E���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�|�!�0�w�}�W���Y���
��1�A܊�
�
�0�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���_��h_�C���d�6�d�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���9�
�
�m�a�8�F���Y����A��B1�Eߊ�g�_�u�u�z�}����H����V9��@����2�u�'�6�$�s�Z�ԜY�Ơ�lS��Z�����"�d�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ѓ�@��GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����Q��D��C���|�!�0�u�w�}�W���Y����G9��V�*���
�0�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ơ�lS��Z�����"�d�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʹ�
�
�c�`�2�m��������[��Z��E���
�g�e�%��}�W�������V�=N��U���`�`�l�
������
���F��G1�*���
�`�b�g�z�l��������lǻN��Xʹ�
�
�c�`�2�m�������]F��X�����x�u�u�9���A����֓�VV��D�����:�u�u�'�4�.�_�������C9��P1������&�f�
�$��N�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�g�;���P����[��=N��U���u�u�u�!�b�h�Nځ�&ù��F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�9�
��k�B���I����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����G9��X�*���
�0�u�&�>�3�������KǻN�����`�l�
�
��8�(�������A	��N�����&�4�
�0�w�-��������`2��C\�����g�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��G݊�&�
�c�|�w�5��ԜY���F�N��*ߊ�c�`�0�e�4�l�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���@���l�
�
�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�!�b�h�Nځ�&ù��Z�=N��U���u�9�9�
�8�����K����9��P1�L���=�;�}�0��0�D؁�&����Q��^��H��r�u�9�0�]�}�W���Y����G��1�����d�`�%�n�]�}�W������P��h��*���u�&�<�;�'�2����Y��ƹF��C1��@��
�
�
�0��.����	����	F��X��´�
�0�u�%�$�:����&����GT��Q��G���u�u�7�2�9�}�W���Yӏ��N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����g�|�|�u�?�3�}���Y���F�[��*��`�0�e�"�f�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��C1��@��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�!�`�b�d�(���&����V��R�����a�
� �g�g��F��T����\��XN�N���u�9�
�
�a�h��������@��S�����f�'�2�g�`�u�W���Y����G	�UװU���x�u�!�`�b�d�(���&����R��P �����&�{�x�_�w�}����L����V9��T�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�m����K��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�D߁�
����O�C��U���u�u�u�u�w�1�(ځ�O�ӓ�lW��R^��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�)�B��@ƹ��9��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�[��*��`�0�d�6�f�<����Y����V��C�U���9�
�
�c�b�8�F���H����Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�c�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�b�3�8�e�t�^Ϫ���ƹF�N��U���!�`�`�l���(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʹ�
�
�c�`�2�l���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�1�(ځ�O�ӓ�lW��N�U���-� �,� ��j����K����9l�N�U���`�`�l�
������
������T��[���_�u�u�!�b�h�Nځ�&¹��9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�b�3�:�o�^���Yӄ��ZǻN��U���3�}�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�`�;���P���G��d��U���u�u�u�9���A����ד�VW�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�!�b�h�Nځ�&¹��F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����lS��1��G���1�0�&�u�j�)���&����V��G_��U���u�:�;�:�g�f�W�������P��h��*���'�&�d�i�w�0�(�������Q��N�Dʱ�"�!�u�|�]�}�W��Y����lS��1��G���e�4�&�2�w�/����W���F�[��*��`�0�g�6�g�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C]�����g�|�|�!�2�}�W���Y���F��C1��@��
�
�
�0�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h[��C���0�g�6�e�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�9���A����ԓ�VW��D��ʥ�:�0�&�u�z�}�Wϲ�&ƹ��
S��h\��ۊ�&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�E؁�
����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���N����lT��G�����_�u�u�u�w�}�W���L����9��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����l��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��C1��@��
�
�
�d�k�}����7����V��V��*؊�0�
�b�a�]�}�W��Y����lS��1��G���d�4�&�2�w�/����W���F�[��*��`�0�g�"�f�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�c�|�|�#�8�W���Y���F���@���l�
�
�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�[��*��`�0�g�"�f�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�;�!�?�l����N�ӓ�F�L�U���;�}�:�
�����H����[��G1�����9�m��|�2�.�W��B�����[��*���d�c�
�g�k�}�G������_	��a1�����c�b�%�u�w�-��������l �������w�_�u�u�8�1�܁����� 9��R��W���"�0�u�9�4��E���&����l��
N��*���&�
�#�
��}����[����F�Y����� �g�l�
�e�a�W��Y����N��T1�����l�`�%�u�w�-��������l �������w�_�u�u�8�/�ށ�����9��R��W���"�0�u�9�4��@���&����l��
N��*���&�
�#�f�g�}����[����F�Y�����3�
�b�l�'�}�J���[ӑ��]F��X��*ߊ� �d�m�
�f�`��������_��h^�����u�e�n�u�w�3����J����Q��h�I���d�u�=�;��2�(���&����S��G_��U���6�;�!�9�e��^ϻ�
���]ǻN��*��d�d�<�3��m�D���Y���F�N�����:�&�
�#�d�m� ���Yے��lW��Q��E���%�}�|�h�p�z�W������F�N�����d�3�
�l�b�-�L���YӖ��V��C1�*���g�a�
�`�k�}����7����#��E��G���
�l�d�%��l��������F�C��GҊ�
� �g�a��n�L���YӖ��V��C1�����l�d�%�u�j�u��������EW��N������3�
�l�b�-�^�ԜY�Ƽ�e��hY�� ��f�
�d�i�w��$���:����lS��Q��C���%�n�u�u�'��݁�&����Q��G_��Hʷ�3�`�d�g���(��s���C9��[\��*���d�e�
�d�k�}����&����l��h����u�=�!�%�>�;�(��A����[�N��U���6�
�!��%�����J����l��h\�Eʢ�0�u�!�%�c�����N���F�_��U���0�_�u�u�w�}�$���5����F��X�� ��`�
�f�_�w�}����&����Z9��D�����3�
�l�`�'�}�J�ԜY���F��h�����#�`�`�e� �8�WǪ�	�Փ�l��h��D��
�g�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�d��m�L���YӔ��l��h�� ��f�
�f�i�w�}�W���YӇ��P	��C1��Dߊ�e�e�"�0�w�)��������l ��W�*��e�u�u�d�~�8����Y���F��G1�����9�d�
�a�g�W�W�������CW��^1��*��b�%�u�h��0�F���&����l��X�����c�1�8�'�6��(���H����CT�=N��U���
�8�d�
��2�(���H����CT�
N�����8�d�
�
�"�l�C؁�KӞ����T�����d�d�n�u�w�.����	�ԓ�l ��_�*��i�u�u�u�w�}��������l*��G1�*���
�0�
�b�g�*����
����^��h�����b�l�e�u�w�l�^ϻ�
��ƹF�N�����%�<�'�2�e�m�L���Yӕ��l��V��*���:�2�;�3��e�D���Y���G��]�� ��m�
�g�:�w�8�(���H¹��U��Z�����_�u�u�0��0�Fׁ�&����S��G\��H���0�
�8�d����������F9��]��Gʭ�'�4�
�:�$��ށ�P���F��[1�����<�3�
�m�b�-�W��Q���� Q��B1�D݊�g�-�'�4��2����¹��l�N�����%�
�
� �f�k�(��E����^��h��*���d�d�
�g�/�/��������_��G�U���&�9�!�%�g�4����A�ד�F�F�����%�m�<�3��e�N���Y����@��C��L���3�
�m�`�'�t�}���Y����G��1�����d�l�%�u�j�W�W���Y�Ư�l
��q��9���
�f�0�e�%�:�E��Y����N��[1�����<�'�2�g�d�u�^��^���V
��d��U���u�&�9�!�'�o����&����l��=N��U���
�8�g�
��(�F��&���F��Z��F���
�b�b�%�w�3�W���&����9��Y�����m�b�%�|�]�}�W���&����
9��Q��M���%�u�h�}�:��C���&����l��V �����!�%�m�<�1��O���	����F�D�����
�
� �d�a��E��Yے��lS��h��*���d�f�
�g�6�9��������Z9��h_�D���|�_�u�u�2����&����lT��1��U��_�u�u�u�w�1��������\��1��E���2�g�l�u�?�3�_���&����
9��E��G��}�|�h�r�p�}����s���F�D�����d�<�3�
�f�d���Y����V
��Z�*��� �d�l�
�e�a�WǪ�	����U��_�����;�u�0�
�:�l�(�������
9��UךU���0�
�8�a�����Kƹ��Z�=N��U���u�%�6�;�#�1�D݁�?����V��_��]���
�8�d�
��8�(��@���F�G�����_�u�u�u�w�����H����lT��B1�Gڊ�f�_�u�u�2����&����lT��1��U��_�u�u�u�w�����H����lW��B1�Dފ�f�"�0�u�$�1����I����V�� ]�E���u�d�|�0�$�}�W���Y����V
��Z�*��� �g�g�
�d�W�W�������CS��^1��*��l�%�u�h�]�}�W���Y����G9��E1�����l�0�e�'�0�o�N������@��C��L���'�2�g�a��t�J���^�Ʃ�@�N��U���&�9�!�%�g�4����H�ԓ� ]ǻN�����8�c�<�3��m�B���Y���D��_��]���-� ��;�"��C���&����C��B1�Bي�f�h�4�
�8�.�(���L����O��[��W���_�u�u�0��0�@�������W��N�U��u�=�;�}��%�"�������R��Y1��!���
� �d�b��n�JϿ�&����G9��[��E���0�&�u�e�l�}�Wϭ�����9��Q��E���%�u�h�}�2���������V��h����0�
�8�b�>�;�(��H����l�N�����%�<�3�
�n�n����D���F�N�����<�<�3�
�n�l�������G��^1�����
�l�l�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�B��I���F��G_�� ��a�
�g�i�w�)���&����A��h�� ��e�
�g�:�w�0�(�������T��^1��*��l�%�|�_�w�}����@����V��h�I���!�%�<�3��d�B���Y����^�� 1�����e�d�%�|�]�}�W���&¹��lT��1��U��_�u�u�u�w�-��������l ��@��U¡�%�<�3�
�n�h����P���A�R��U���u�u�u�4��2����˹��9F���*ۊ�
�d�<�3��k�@���Y���D��_��]���
�
�
� �f�e�(��DӇ��P	��C1��Gي�|�0�&�u�f�f�W�������l��1�����b�f�%�u�j��Uϩ�����\��hY�� ��g�
�d�h�6�����&����lV�R��U��n�u�u�!�'�l��������P��h�I���e�u�=�;��2�(���&����S��G_��U���6�;�!�9�e��^ϻ�
���]ǻN�����e�3�
�`�o�-�W��Q����]	��h����b�<�'�2�f�i�W���Y����\��h��*���_�u�u�8��l����L�ғ�F���*���<�
�0�!�%�/����Q����T����*���3�
�`�m�'�t�A���B�����h\�����c�d�%�u�j�.��������V��EF�����}�;�<�;�3�4�(���&����J��G�U���!�%�g�
�"�l�E߁�H���@��[�����6�:�}�0�>�8��������Z*��^1�����:�
�
�0��i�E��M����F�C��Gފ� �g�f�
�d�a�W���Y�����h_�� ��g�
�f�"�2�}����Hʹ��lT�� 1��]���h�r�r�u�;�8�}���Y���G��_�� ��g�
�d�_�w�}����L����V��h�I���!�%�f�<�>�4����@�ӓ�F�� �����3�
�e�d�'�t�}���Y����Q��B1�Eي�g�i�u�!�'�o�(���K����CT��Y
����� �d�d�
�e�f�W�������9��Q��E���%�u�h�w�u�*����
����WN��h��9����!�m�
�9�8����H����_��h�U���<�;�1�4��2�����ޓ�O��[��W���_�u�u�8��e����N�ѓ�F�F�����d�3�
�b�f�-�W�������@W��B1�Aߊ�g�n�u�u�#�-�Eׁ�&����R��G]��H���8�
�a�3��m�D���Y�Ƽ�W��h_��*���g�d�
�f�l�}�WϪ�	����U�� Y�����h�}�:�'�$����Oʹ��	��Y�����3�
�b�f�'�t�}���Y���� V��B1�Mۊ�g�i�u�!�'�o�(���H����CT��Y
�����l�3�
�b�b�-�^�ԜY�Ƹ�C9��h��G��
�d�i�u��%�"�������R��Y1�����d�3�
�l�n�-�_���Y�ƨ�D��^����u�8�
�f�1��@���	���N��G1�*���d�m�
�g�6�9��������_��G�U���!�%�f�
�"�l�Gځ�K�����E��*���d�l�
�g�8�}����
����lW��1��\�ߊu�u�8�
�b�;�(��H����[�C��Fފ� �d�e�
�e�<�Ϫ�	����U�� [�����_�u�u�8��k��������Z9��h_�B���u�h�}�8���F�������S��N��ʡ�%�d�<�<�>�;�(��H����l�N����
� �d�g��-����E�ƭ�l��D��ߊ�n�u�u�!�'�n�(���H����CT�
N�����`�3�
�m�f�-�W���Y���� P��B1�Gߊ�g�n�u�u�#�-�Dׁ�����R��h��D��
�g�i�u�#�-����&����lW��1��U���u�8�
�
��l����&����l��d��Uʡ�%�f�<�<�>�;�(��L����[�L�����}�:�
�
��(�F��&�����T�����g�
�|�0�$�}�G��Y����^��1�����4�
�
� �f�n�(��E����^��h�����
�b�b�%�w�3�W���&¹��ZT��h��D��
�g�n�u�w�)���&����V��G_��Hʦ�1�9�2�6�!�>����������^	��¼�
�0�
�a�d�q�C���s���G��_�� ��d�
�d�i�w�)�(�������P������� �&�2�0��n����H����P��UךU���8�
�g�3��e�D���Y���G��Z�� ��e�
�g�4�3�)���&����Q��G\����u�8�
�f�1��B�������VF������!�9�`�g�]�}�W���&�ғ�F9��W��G��u�!�%�a��(�F��&����]��Z��F���
�`�e�%�~�W�W�������l ��_�*��i�u�!�%�c�����N����]��E�� ��d�
�g�n�w�}����MĹ��lW��1�����u�h�4�
�8�.�(���&��ƹF��Z��M���
�m�`�%�w�`�_���&�ӓ�F9��_��Gʴ�1�!�%�a��(�F��&���9F���*ߊ�
�
�
� �f�n�(��E���F��R ������3�
�l�b�-�W���	����@��AV��3���9�0�w�w�]�}�W���&����S��G_��Hʦ�1�9�2�6�!�>����������^	��¼�'�2�d�f�~�k�^��Y����^��h��D��
�g�i�u�f�}����Q����V��d1�� ���;� �
�a�>�����&¹��lW��1��\��&�2�0�}�'�>��������u#������w�_�u�u�:��(�������P��h�I���d�u�=�;��2�(���&����R��GZ��U���6�;�!�9�o��^ϻ�
���]ǻN�����
�g�<�3��k�F���Y���D��_��]���
�
�
� �f�j�(��DӇ��P	��C1��M���|�0�&�u�g�f�W�������l��^1��*��b�%�u�h�u�� ���Yۊ��l0��h��D��
�a�h�4��2����˹��F��D��E��u�u�!�%�>�4����&����l��S��D���=�;�}�:�����Iƹ��[��G1�����9�m�e�u�;�8�U���s���G��D1��*���f�%�u�h�$�9��������G	��E�����;�<�;�1�6�/����&����lT��h�����a�l�y�a�~�W��������9