-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�?����P��1��@���3�`�f�`�2�m������ƹF��R �����u�u�u�u�w�}��������F������o�u�7�:�<�f�}���Y���F�S�����u�u�u�;�2�8�W��J���F�N��U���4�<�!�u�w�}�W�������	[�NךU���u�u�u�u�2�����Y����Z��P��O���_�u�u�n�]�}�W�����ƹF�N��U���'�u�u�u�w�3��������l��C�����!�x�u�:�9�2�G��s���F�N��E���u�u�o�<�w�)�(������F�N��Uʤ�u�u�u�u�m�2�ϭ�����Z��R��±�<�!�x�u�8�3���B���F�N�����u�u�u�u�9�.��������V��EF�����x�u�:�;�8�m�L�ԜY���F�T�U���u�o�<�u�#�����B���F�N�����u�u�u�o�>�}��������E��X�����=�d�1�"�#�}�^���Y���F���U���u�u�u�;�$�9������ƹF�N��U���u�u�u�u�m�4�W���&����PFǻN��N���;�u�;�<�.�}�}������P��RN��ʺ�u��c�e�f�;�G���L����lS��[��*ڊ�4�u�&�_�$�:��������G��N�����2�6�#�6�8�u� �������\��XN�N���,�0�8�8�6�/�Ϸ�Y����JF������&�/�x�|�8�}��������E��X�����!�x�u�:�9�2�G��s����V��V�����'�8�o�8�:�<����s����A��C�����4�&�,�0�m�.����B���G��B�����'�8�!�9�w�;����CӐ��Z��RN��Uȷ�:�>�'�8�l�<��������R��C��U���!�<�2�_�#�/����Y����@��RN��U���u�u�4�<�5�8��������C��V�����0�� ����(���0����l4��x8��U���!�<�2�_�5�:��Զs����A��T�����4�1�e�u�%�>��������F��R	�����u�u�1�'��0�W������l�D�����&�!�4�&�6�8����Y�����-��#������4�3�m�W�������I�N���ߊu�u�u�u�w�<�������F��C����u�e�|�_�w�}�W������F�N��U���'�
�8�u�j�<���s���F��SN��N���&�;�=�&�$�)��������]l��SN�����&�_�%�8�:�/�(�������	F��X�����9�|�u�7�0�3�}���Y���P
��R��ʴ�1�6�>�h�p�z�W������F���]���u�u�d�|�#�8�W���Y���F��I���4�}����	�0�������l��G����u�u�u�;�w�;�}���Y����Z ��R �����0�&�_�_��8��������@9�������u�6�>�u�]�8����Y����UF��[�����u�;�u�9�w�}�F�������F�N�����6�d�h�r�p�}����s���F�N�����"�d�h�r�p�}����s���F�N��U���'�8�����2���Q����O�S��D���u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}�����Ƽ�\��DUװ���u�!�n�_��?����0����9��'��0Ħ�1�9�2�6�f�k�Y���B���G����C���d�3�e�3�b�?����J�ӓ�lV��Dd��Uʲ�;�'�6�}�w�}�W���=����Z��T��;����u�h�f�l�}�W���Yӧ��A��e��������m�}�L���Y���'��E��"���=�o�����M���P���F��E�����u�u�u�0�2�}�W���*����|!��d��U���u�6�>�o��}�#���6����9F�N��U���'�&�e�o��}�#���6����e#��x<�����&��1�=�z�l�3���-����l�N��Uʶ�e�o��u���8���B���F��Oʚ�������!���6�Έ�G��S��X�����u�~�W�W���Y�ƭ�W��D_��U���������4���Q����V��^
��U���u����g�f�W���Y����VW�'��&������_�w�}�W�������z(��c*��:���n�u�u�u�w�9�W���7ӵ��l*��~-��0�����!��3�5�Z��=����|F��U�����;�<�,�_�6�>��������R�������a��c�
���(���&ƹ��9��N�����u�:�%�;�9�}�6��I����lV��h[�� ���
�e�
�
��<�W���Y���F��X��]���u�u�u�u�w�>���0�Ɵ�w9��p'�����u�u�u�u�w�9����Y����g"��x)��*�����_�u�w�}�W���Y����	F��=��*����n�u�u�w�}�W�������|3��d:��9�������l�}�W���Y�����E_��U���������4���B���F�N��U���u�u�����0���s���F�N�����u������4���:����9F�N��U���u�0�u�u���3���>���9F���U���%�;�;�n�]�W����s���^'��^��C���
�
�
� ���Gځ�&ù��^9��N�����;�;�u��a�m�Fٸ�I����l��h[��Eߊ�
�
�4�_�w�}�������9F�N��U���u�k�6�>�]�}�W���Y����F������e�_�u�u�w�}����GӅ��l�N��Uʤ�u�k�$�y�w�}�W�������[�V
�����y�u�u�u�w�>�F��Y����9F�N��U��h�u�d�_�w�}�W��������Uװ���4�6�<�0�#�/�L�Զ