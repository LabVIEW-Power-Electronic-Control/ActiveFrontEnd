-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�8����_��1��F���3�f�d�m��<�W���s���T��E�����u�u�u�u�w�8�(������	F��E��U��w�9�6�w�w�}�W���Y�����S��U���o�<�!�2�%�g�W��Y���F�N��U���1�=�u�u�m�4�������]�N��U���u�u�8�8�$�'�W���Cӏ��V��T��G���u�|�u�u�w�-����s���F�N����u�u�o�<�w�)�(�������P�������d�1�"�!�w�t�W���Y���F��R^��U���u�u�;�&�3�1����Y���F�N��E���u�u�u�u�"�}��������E��X�����=�d�1�"�#�}�^�ԜY���F�V
��D���u�o�<�u�#�����&����\��@����1�"�!�u�~�}�W���Y�����N��U���u�;�&�1�;�:����Y���F�
�U���u�u�u�;�$�9��������G	��S�����u�:�;�:�g�f�}���Y���F��N��U���o�<�u�!��2���s���F�N��U���u�u�o�:�#�.��������V��EF�����x�u�:�;�8�m�L���Y���F��[��U���u�o�<�u�#�����Y���O��=��U���<�,�u�_�6�>��������A��X��E��`�d�3�e�1�n����J����9��ZN��U���<�;�9�4�3�m����Cӕ��l
��^�����'�4�<�!�z�}�������l��P ��U���'�
�8�u�w�)�(�������P�������d�1�"�!�w�t�W��	�ơ�^9��E�����'�4�u�e�#�}�������F����*���<�
�0�!�%�u� �������\��XN�N���=�'�1�#�%�<��������^��V���ߠ4�!�<� �2�.��������VF��D����_�!�'�7�#�}��������_��QN����#�'�4�9�w�.�U�������^D��V�����0�'�8�&�.�8�Mϭ�����9��E�����4�
�!�9�w�;����CӐ��Z��RN��U���
�,�0�_�#�/����Y����e'��y:��0���������Mϭ�����9l��P�����0�:�,�4�4�.�(���������T��U´�1�e�u�7�0�3�W���YӇ��AV��Z��Hʴ�1�e�_�x�.�)����Y����@
��R1�����u�u�<�u���(���<����R��G��U���
�<�0�d�w�5����Y���F�V
��E���%�i�u�:�?�/�W���^���9F�N�����_�u�u�u�w�}����I����Z�V
��E�ߊu�u�u�;�w�;�}��� ����@��C�����0�:�_�;�w�/����B���^��E�����&�e�u�'�4�.�Wǽ����Q��YNךU���3�}�9�r�!�3�W���Y����F�G�����u�u�u�u�>�}���D����F��R ��U���u�u�u�u�&�}�JϬ�ۥ��e9��c+��'´�1�e�!�%�~�}�W���Y����]��QUךU���;�u�3�_�9�}����
��Ɠ^��E�����&�2�4�1�f�}����
����W��N�����_�u�u�u�3�/�(���Y����W��d����=�&�&�!�6�.������ƹF���]��������<���Y�ơ�^9��M��\ʡ�0�_�u�u�w�}�WϿ��ד�^�
N�����&�h�u�e�~�W�W���Y����l�N��U���u�1�'�
�:�}�JϿ�����F�N��ʼ�n�x�&�;�?�.�Ϫ�����G��Yd��ʥ�:�0�&�_�'�0����&����@��N�����&�}�9�|�w�?����s���Z �T�����!�4�1�6�<�`�P���Y����9F�N��U���}�0�u�u�f�t����Y���F�N��U���}�0�u�u�f�t����Y���F�N��U���u�4�}����#���+ۇ��AW��Z��U��1�n�_�u�w�}�W���Y����Z ��N��U���u�u�$�u�j�/�ǝ�7����g#��eF�����!�%�|�u�w�}�W�������U]ǻN�����3�_�;�u�%�>���s������dװ9���4�,���l�(�ϗ�<�ȿ�W9��P��D��{�9�n�_�9�4�ϳ�8����_��1��F���3�f�d�m�w�.�W�������Z�=N��U���u�4�4�<�#�}�W���<����	[�UךU���u�u�1�'�$�����Cӯ��v!��T��G�ߊu�u�u�u�3�/�������/��r)��U��d�n�u�u�'�/�W�ԜY���F��D��Oʜ�u��
���f�W���Y����_�'��&������_�w�}�W�������@V�'��&���������_�������Z��C��U�����e�n�w�}�W������/��d:��9����_�u�u�w�}�G��6����g"��x)��*������!� �9���HӢ��}2��G�U���u�u�4�1�2�.�W���7ӵ��l*��~-��0�����1�0�$�4����Y�ƈ�d(��^����u�u�u�0�w�}�9ύ�=����z%��N��U���"�d�o��w�	�(���0��ƹF�N��D���u��
���(���-����R��^
��U���u����g�f�W���Y����F��x;��&���������_�������[F�N��"���u�|�n�0�3�8����B���P��R�����'�=�:�u�g�k�B���֓�lU��B��*��a�<�_�u�w�2�����ơ�rP��_��*ڊ�
�
� �
��e�C���ӏ��F�N�����u�_�u�u�w�}�W�������z(��c*��:���n�u�u�u�w�}�WϿ����/��d:��9�������l�}�W���Y�����T��;ʆ�����]�}�W���Y���BV�!��U���
���
��	�%�ԜY���F�N����o��u����>���<����l�N��U���u�6�d�o��}�#���6����9F�N��U���u�d�o��w�	�(���0����p2��d��U���u�u�u�"�f�g�>���-����t/��=N��U���u�u�u�d�m��#ύ�=����z%��r-��'��u�u�0�1�4�0������Ɠ9��^ ךU���e�c�`�d�1�m��������lW��1�����o�u�:�%�9�3�W���O����
 ��h��*���
�
�m�a�%�0�W���	����^��d��U���u�6�>�h�w�1�[���Y�����E^��Kʴ�1�0�&�y�w�}�W������F��BךU���u�u�e�h�w�m�}���Y���R��N��U���'�&�d�_�w�}�W��������d��U���u�1�u�k�3�q�W���Y����VW�	N��D�ߊu�u�u�u�f�`�W��B���WF��T�����'�n�_�