-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�8����_��1��F���3�f�f�`�2�m������ƹF��R �����u�u�u�u�w�}��������F������o�u�7�:�<�f�}���Y���F�S�����u�u�u�;�2�8�W��J���F�N��U���4�<�!�u�w�}�W�������	[�NךU���u�u�u�u�2�����Y����Z��P��O���_�u�u�n�]�}�W�����ƹF�N��U���'�u�u�u�w�3��������l��C�����!�x�u�:�9�2�G��s���F�N��E���u�u�o�<�w�)�(������F�N��Uʤ�u�u�u�u�m�2�ϭ�����Z��R��±�<�!�x�u�8�3���B���F�N�����u�u�u�u�9�.��������V��EF�����x�u�:�;�8�m�L�ԜY���F�T�U���u�o�<�u�#�����B���F�N�����u�u�u�o�>�}��������E��X�����=�d�1�"�#�}�^���Y���F���U���u�u�u�;�$�9������ƹF�N��U��u�u�u�u�w�(�W���&����P9��T��]���1�=�d�1� �)�W���s���F�N�����u�u�u�u�9�.�������F�U�����0�!�!�n�]�W��������A��C��ʸ��b�d�l���(܁����� V��R1�����<�u�_�<�9�1����I����\��C
�����
�0�!�'�6�4���Y����G	�U�����4�u�1�'��0�W�������T��A�����"�1�=�d�3�*����P����J��Z�����,�<�u�'�6�}�GϪ�Y����@��_�����!�
�:�<��8����Q����G�
�����e�n�_�=�%�9��������A��N�����'�,�_�4�#�4����
����R��N��Oʦ�'�;�n�_�#�/����Y����A��C��U���'�8�o�#�%�<����
�Į�\��E��N��!�<� �0�%�0��������G��PU�����7�!�u�4��)����Ӕ��\��V�����<�u�0�
�.�8�}�������VF��b'��9���
������:���5����G��PUװ���;�_�_�0�8�$����
����R��T�����&�u�4�1�g�}�������F��S
��*���u�h�4�1�g�W�Z�������@F��V �����:�3�u�u�w�4�Wǝ�7����g#��eF����u�u�0�
�>�8�F�����ƹF�N��Uʴ�1�e�!�%�k�}�������A��UךU���u�9�0�_�w�}�W���YӇ��AV��Z��Hʴ�1�e�_�u�w�}�������@��_��ʡ�4�&�4�0�8�W��������@]ǑG1�����
�6�0�&�g�}����
����_�d�����_�u�u�3��1�P����ƭ�WF��\N��R��u�=�;�u�w�}�WϷ�Yۅ��[�I�����u�u�u�u�w�}�Wϯ�Y����R��x ��<�����4�1�g�)����Y���F���U���_�u�u�;�w�;�}���Y����V��=d�����
�6�0�&�0�<���Y����V�������_�0�<�_�w�}�W���¹��CF�����x�&�;�=�$�.����
����l	��=N��U���3�}����	�0�������F�Z�����x�|�!�0�]�}�W���Y����W��h��U��}�!�0�&�j�}�G���s���F��D��U���u�u�u�u�3�/�(���Y����W��d��U���0�1�<�n�z�.����
����A��[��*���0�1�%�:�2�.�}������J9��T��*��%�:�0�&��1�^�������l�N��U¶�>�0�0�!�6�9����D����F��R ךU���u�u�3�}�2�}�W��PӒ��]FǻN��U���u�u�3�}�2�}�W��PӒ��]FǻN��U���u�u�u�u�6�u�8���0����v4��S
��*���|�u�h�1�l�W�W���Y���F��SN��N���u�u�u�u�w�,�W������|(��~ ��2���4�1�d�!�'�t�W���Y����������u�;�u�3�]�3�W�������9l��Y
����_��7�4�.��2������v#��D�����6�d�c�{�;�f�}�������'��_����3�f�7�3�d�n�B���Iӏ��F�P�����}�u�u�u�w��������/��r)��U��f�n�u�u�w�}�6�������]��N��!����o�u�n�w�}�W���8����@��S��Oʜ����o�w�t�}���Y����NǻN��U���0�0�u�u���3���>����F�N�����o��u����>��Y���F��S
����o��u����>���<����'��E��"���=�x�d�� �	�W���s���F�T�Oʜ�u��
���f�W���Y����F��x;��&���������_�������[F�N��"���u�|�_�u�w�}�W�������\��yN��1��������u����
����G�_��:����e�n�u�w�}�WϽ�H����}F��s1��2���_�u�u�u�w�8�W���7ӵ��l*��~-�U���u�u�1�u�w��$���5����l0��c!��1����1�=�x�f�� ���Y����F�N�����u� �u����>���<����"��V9�����u�u����m�^����Ʃ�G��d�����!�6� �0�6�>�W���ç��W��Q1�����7�3�f�f�b�8�GϷ�s���P	��X ��ʸ��b�d�l���(܁����� V��R1�����<�_�u�u�w�}����Q���F�N��U���u�u�����0���s���F�N�����e�o��u���8���&����|4��N��U���u�u�6�e�m��W���&����p]ǻN��U���u�u�e�o��	�$���5����l0��c!�����u�u�u�u�w�9����Y����g"��x)��*�����_�u�w�}�W���Y����	F��=��*����n�u�u�w�}�W�������z(��c*��:���
����]�}�W���Y���D��N��U���
���n�w�}�W���Y����F��x;��&���������^�ԜY�Ʃ�WF��Z�����_�_�7�2�9�}�Wϳ�8����_��1��F���3�f�f�`�2�m����,���P	��X ��ʸ��b�d�l���(܁����� V��R1�����u�u�%�'�w�<�W�ԜY���F��\N��U���y�u�u�u�w�<���D�ƭ�W��D^�U���u�u�6�e�j�}���Y���F��N��U��_�u�u�u�w�9����GӇ��A��BךU���u�u�0�u�i�>�F�ԜY���F��S����u�u�u�u� �l�J�����ƹF�N��D��u�d�n�_�9�}��������A��=d