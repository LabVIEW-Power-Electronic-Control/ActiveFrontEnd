-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��G���Jˀ��l ��U1����g�&�f�
��(����	ӏ��F�P�����}�u�u�u�w��W���Y���	F��C����u�a�_�u�w�}�W���&����vF������u�h�f�_�w�}�W����֓�z"��T�����0�u�h�f�l�}�W���Yӂ��9��s:��Oʼ�!�2�'�o�w�o�}���Y���W	��h9��!���u�;�0�0�w�`�D�ԜY���9F������u�u�u�u�4�6�W������G��X	��N���u�u�u�'�$�)�MϷ�Yӕ��l
��^�U���u�u�6�u�w�g����
����\��d��U���u�1�;�u�m�4�Wϭ�����Z��R��±�;�
���z�}�������9F�N��U���d�u�u�;�w�)�(�������P��
��D�����d�1� �)�W���s���F�S��U��:�!�&�1�;�:��������W	��h9��!���u�:�;�:�g�W�W���B������^����6�<�0�!�%�}�����ơ�V��v]��*ڊ�&�7�f�;��o���&����_
��D�����u�x�x�x�z�p�Z��T���K��X�����u�x�x�x�z�p�Z��T���l�N�����0�!�8�a�a��O���&����@��1�����&�
�g�<�]�}�W���Y����NǻN��U���u�u�6�>�w�}�W���Y���F���U���
�:�<�n�w�}�W���Y����P
��YN��U���u�u�u�u�m�4�Wϭ�����Z��N��U���u�u�&�4�>��(������F�N��Uʦ�1�9�2�6�]�}�W���Y���@9��^��*���!�u�u�u�w�}��������T��A�����d�1�"�!�w�t�}���Y���F�D1�����
�#�9�1�w�}�W����ƿ�W9��P�����u�u�u�u�w���������G�N��U���;�u�!�
�8�4�(������F��@ ��U���_�u�u�u�w�}�W�������V��C1�����u�u� �u�#�����B���F�N��U���-�&�'�&�;�����Y����F��C
�����
�0�!�'�d�}�������F�N��\�ߊu�u�;�u�8�-����B���K�C�X���x�x�x�x�z�}����Y����R
�C�X���x�x�x�x�z�}�Wϭ�����R��N��U��&�1�9�2�4�W�W���������\��U���u�!�
�:�>�f�W���
����_F��C�����o�&�1�9�0�>�}���Y����R
��h�����u�u�!�
�8�4�(������F��@ ��U���_�u�u�<�9�1��������\��C
�����n�u�u�&�0�<�W�������F��D�����6�#�6�:��l��������l�N�����u�
�#�9�3�}�W���&����P]ǻN�����9�'�!�4�6�}�Mϭ�����Z��R����u�:�;�:�g�f�W���
����_F��Y^�� ��o�&�1�9�0�>�����Ψ�]V��~*��X���:�;�:�e�l�}�Wϭ�����W��h��D��&�1�9�2�4�+����Q����l1��c&��U���;�:�e�n�5�:����Y���K�C�X���x�x�x�u�9�)��������K�C�X���x�x�x�u�w�0�C��8�ު�9��h�����3�9�
�&��o�������]����E���f�3�e�4��.��������W��\ךU���:�!�8�%��}�W���YӇ��XF�N��U���u�u�u�h�w�>��ԜY���F��[��U���u�u�u�u�w�}�IϿ�����9F�N��U���-�&�4�!�6�4�W���Y���R9��V��Y���u�u�u�&�6�4�(�������F�N��U���1�!�y�u�w�}�Wϭ�����Q9��V��U���u�h�u�
�!�1��ԜY���F��V��*���1�!�u�u�w�}�Iϼ�����l�N��Uʸ�4�<�
�0�"�)���������A���ߊu�u�u�u��%����
����G��VN��Kʧ�!�4�4�u�w�t�}���Y���K�C�X���x�x�x�u�$�4�������K�C�X���x�x�x�u�w�<����Y�����d��Uʴ�9�0�u�u�j�>�L���YӇ��E��SN�U��n�u�u�4�#�<����D�Ψ�]V��~*��X���:�;�:�e�j�}�G�������N��Y^�� ��h�}�1�;���#��Y����G	�S�R��|�u�'�}�>�m����Y���W��h9��!���u�:�;�:�g�`�Wȋ�P����_��S��*���d�_�u�u��+����E���]ǻN��*���!�u�i�u�3�3�(���-����W	��C��U��r�r�u�=�9�u����&����[�
��D�����d�1� �)�W���G����O�X�����
� �d�h��9�ށ�0����F��@ ��U���k�r�r�|�w�1�Ϻ�¹��UW��N�����u�u�u�h�%�)����s���K�C�X���x�x�x�x�z�}����Y����V�C�X���x�x�x�x�z�}�WϮ�����N��\G�����_�u�u�u�w�;������������U���d�u�=�;�w�}�W���Y����UF��S��D���=�;�u�u�w�}�W���Y����Z��U��U��1�;�n�u�w�}�W���Y�����1�����h�1�;�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���4�6�<�0�#�/�L�