-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�?����P��1��@���3�`�g�f���(���Y���F�P�����_�u�u�u�w�}�W���&����F�N�����u�h�w�9�4��W���Y���F�
�����u�u�o�<�#�:���Y���F�N��U���4�<�!�u�w�}�W�������	[�NךU���u�u�u�u�2�����Y����Z��P��O���_�u�u�n�]�}�W�����ƹF�N��U���'�u�u�u�w�3��������l��C�����!�x�u�:�9�2�G��s���F�N��E���u�u�o�<�w�)�(������F�N��Uʤ�u�u�u�u�m�2�ϭ�����Z��R��±�<�!�x�u�8�3���B���F�N�����u�u�u�u�9�.��������V��EF�����x�u�:�;�8�m�L�ԜY���F�T�U���u�o�<�u�#�����B���F�N�����u�u�u�o�>�}��������E��X�����=�d�1�"�#�}�^���Y���F���U���u�u�u�;�$�9������ƹF�N��U���u�u�u�u�m�4�W���&����PFǻN��N���;�u�;�<�.�}�}������P��RN��ʺ�u��c�e�f�;�G���L����lS��]�����'�8�<�u�]�4��������l��T�����:�<�
�0�#�/��������W	��C��\���!�%�u�0��/����
Ӈ��R�N��U���
�<�0�d�w�;��������l��C��]���1�=�d�1� �)�W���Y����A��A�����u�4�u�u�2�����B���G��B�����'�8�!�9�w�}��������G��U��U���
�4�&�,�2�2�W���Y�ƺ�A��[�����9�6�
�4�u�W��������A��D����&�'�;�n�6�)����Ӕ��l��[��ʧ�8�o�#�'�6�1�W�������J��=�����!�u�����#���>����a9��z!��9��&�'�;�n�]�8����s����\��V����� �'�
�o�'�2����Q����O�U�����u�u�4�1�g�)���Y����]Ƕ�����<�u�'�;�;�)�(���s���F��F��;������}�3�/�^�������Z��G�����u�u�u�u�w�}����&����[�X�����k�r�r�n�w�}�Wϻ�
��ƹF�N��Uʴ�1�e�!�%�k�}����B���F��Y
���߇x�,�!�0�>�}��������\��Y
�����&�n�_�
�2�2��������\��E�����6�>�u�_�2�4�W���Yӏ���������;�u�9�u�w�l�^Ϫ����F�N��U¶�e�h�r�r�w�5��ԜY���F�N��U��'�8�����2���Q����9��GG�U���u�u�u�0�3�4�L���YӃ����=��U���6�&�n�_�'�0����&����@��N�����&�}�9�|�w�?����s���Z �T�����!�4�1�6�<�`�P���Y����9F�N��U���}�0�u�u�f�t����Y���F�N��U���}�0�u�u�f�t����Y���F�N��U���u�4�}����#���+ۇ��AW�T����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9�������A	��D���1�'�9�_�]�4����Y����l��RN��0���!�
�:�<��l�C�������]��NN��3���c�
�
������&����l����U���2�;�'�6��}�W���YӢ��R1��C��U�����u�h�f�W�W���Y�ƍ�W��D<�����u����w�`�C�ԜY���F��S�����!�u�u����W��K��ƹF��X��]���u�u�u�'�$�)�Mϗ�Y����)��tUךU���u�u�9�u�w��$���5����l�N��Uʴ�1�0�&�u�w��$���5����l0��c!��4���0�&�<�!�w�}�W���7���]ǻN��U���0�u�u����;���:���F�N��U��� �u��
���(���-����R��^
��U���u����g�f�W���Y����W��D�Oʜ�u��
����2���+ۧ��A��`�����d����w�t�}���Y���P��N��U���
���n�w�}�W������/��d:��9����_�u�u�w�}�F��0�Ɵ�w9��p'��#����}�4�4�>�)�W���Y����g)�G����0�!�!�n�]�/����������_N��U���c�e�d�3�g�;�B����ӓ�
U��R1��ߊu�u�:�%�9�3�W���O�֊� ��h��*���
�
�l�d�2�m�������F�N�����_�u�u�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�w�}����I����}F��s1��2������n�w�}�W���Y����VV�'��&������_�w�}�W���Y�ƽ�\��b:��!�����
����}���Y���F�V
��D���u��
���(���-����F�N��U���6�d�o��w�	�(���0��ƹF�N��U���d�o��u���8���&����|4��N��U���u�u�"�d�m��W���&����pO��N�����6�8�:�0�#�W�}����ƹF��v(�E��3�e�3�`�5�;�B��J¹��9��Z1��O���:�%�;�;�w��A���Hŀ��l ��h��*ߊ�l�d�0�e�%�0�W���	����^��d��U���u�6�>�h�w�1�[���Y�����E^��Kʴ�1�0�&�y�w�}�W������F��BךU���u�u�e�h�w�m�}���Y���R��N��U���'�&�d�_�w�}�W��������d��U���u�1�u�k�3�q�W���Y����VW�	N��D��_�;�u�'�?�)������Ɠ