-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�g�e�f���}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e��!�:�$�8�G��6����g"��x)��*�����}�d�3�*����P���F��1�����&�0�e�4��1�W���,�Ɵ�w9��p'�����u�
�
�6�>�3�(���Y�ƃ�gF��s1��2������u�d�}�������9F���*���<�;�
�
��-����Cө��5��h"��<��u�u�%�e��)�������)��=��*����
����u�FϺ�����O��N������!�:�&�2�o��������|3��d:��9����_�u�u���������� F��x;��&���������W��Y����G	�UךU���
�
�6�<�9��(܁�	����\��b:��!�����n�u�w�-�G�������l��T�� ����
�����#���Q����\��XN�N���u�%�e��#�2����M����E
��N��!ʆ�����]�}�W���&����\��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
��>����&����R��[
��U���u��
���f�W���	�֓�P��Y��*���u� �u����>���<����N��
�����e�n�u�u�'�m�6�������lP��G1����������4�ԜY�Ƽ�9��C�����b�o�����;���:����g)��]����!�u�|�_�w�}�(߁�����@9�� 1��*���u�u� �u���8���B�����h/�����
�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�I����Z	��h��*���#�1�o����3���>����F�G1��4���:�&�0�l�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����r��X �����4�
�9�u�w��W���&����p]ǻN��*ي� �%�!�
��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lU��B�����
�
�%�#�3�g�8���*����|!��d��Uʥ�f��!� �$�8�F��6����g"��x)��*�����}�d�3�*����P���F��1�����&�0�d�4��1�W���,�Ɵ�w9��p'�����u�
�
� �'�)�(���Y�ƃ�gF��s1��2������u�d�}�������9F���*���%�!�
�
��-����Cө��5��h"��<��u�u�%�f��)�������)��=��*����
����u�FϺ�����O��N������!� �&�2�n��������|3��d:��9����_�u�u����������F��x;��&���������W��Y����G	�UךU���
�
� �%�#��(ہ�	����\��b:��!�����n�u�w�-�D�������l��T�� ����
�����#���Q����\��XN�N���u�%�f��#�(����L����E
��N��!ʆ�����]�}�W���&����F��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
��(����&����R��[
��U���u��
���f�W���	�Փ�F��C��*���u� �u����>���<����N��
�����e�n�u�u�'�n�8�������lQ��G1����������4�ԜY�Ƽ� 9��C�����m�o�����;���:����g)��]����!�u�|�_�w�}�(܁�����@9��1��*���u�u� �u���8���B�����h!�����
�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�J����C��h��*���#�1�o����3���>����F�G1��:��� �&�0�d�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l)��G��*���e�4�
�9�w�}�"���-����t/��=N��U���
�4� �9�8�)����&����z(��c*��:���n�u�u�4��8�Mϗ�Y����)��tUךU���
�
�4� �;�2����&����R��[
��U��������W�W���&ǹ��]��t�����0�d�o��w�	�(���0����p2��F�U���;�:�e�n�w�}����4����_%��C��*���
�%�#�1�m��W���&����p]ǻN��*ފ�4� �9�:�#�2�(���Y�ƅ�5��h"��<��u�u�%�a��3��������l��h�����o��u����>��Y����lR��V �����!�:�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����~��V�����9�0�f�4��1�W���7ӵ��l*��~-�U���%�a��;�6���������\��yN��1�����_�u�w��(�������]��[1��A���
�9�u�u���3���>����F�G1��8���4��;�'�;�8�B��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����h#�� ���:�!�:�
����������}F��s1��2���_�u�u�
��<��������_9��N�<����
���l�}�WϮ�M����F��X �����
�
�%�#�3�g�>���-����t/��=N��U���
�4� �9�8�)����&����z(��c*��:���
�����l��������l�N��A���;�4��;�%�1��������WF��~ ��!�����n�u�w�-�B�������lV�'��&���������W��Y����G	�UךU���
�
�4�2���(������/��d:��9����_�u�u������&����	F��=��*����
����u�FϺ�����O��N������;�0�0�f�<�(���Y�ƅ�5��h"��<��u�u�%�`��3����K����}F��s1��2������u�d�}�������9F���*���2�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�4�0��(���Y����g"��x)��*�����}�d�3�*����P���F��1�����0�f�4�
�;�}�W���*����|!��d��Uʥ�`��;�0�2�i�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����lS��V ��*���
�%�#�1�m��W���&����p]ǻN��*ߊ�4�2�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����a��R1��@���
�9�u�u���3���>����F�G1��'���0�0�c�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�L����T��hX�����1�o��u���8���B�����h<�����
�u�u����;���:����g)��]����!�u�|�_�w�}�(ځ�����V9��V�����u������4�ԜY�Ƽ�9��Y	����o��u����>���<����N��
�����e�n�u�u�'�h�%�������l��A��Oʜ�u��
���f�W���	�ӓ�R��h��U���������!���6���F��@ ��U���_�u�u�
��<����&ʹ��l��T��;ʆ�����]�}�W���&����^��E��*���u������4���:����U��S�����|�_�u�u����������l��h�����o��u����>��Y����lP��V�����&�0�d�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�O����R��R�����4�
�9�u�w��$���5����l�N��C���'�8�!�'���W���7ӵ��l*��~-��0����}�u�:�9�2�G��Y����lP��V�����&�0�g�4��1�W���7ӵ��l*��~-�U���%�c��'�:�)����&����z(��c*��:���
�����l��������l�N��C���'�8�!�'���(������/��d:��9����_�u�u����������l��T��;ʆ�������8���Iӂ��]��G�U���%�c��'�:�)����&ǹ��l��T��;ʆ�����]�}�W���&����@9��N�<����
�����#���Q����\��XN�N���u�%�b��>�.��������WF��~ ��!�����n�u�w�-�@�������lW�'��&���������W��Y����G	�UךU���
�
�4�;���(������/��d:��9����_�u�u������&����	F��=��*����
����u�FϺ�����O��N������<�&�0�e�<�(���Y�ƅ�5��h"��<��u�u�%�b��4����J����}F��s1��2������u�d�}�������9F���*���;�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�4�9��(���Y����g"��x)��*�����}�d�3�*����P���F�� 1�����0�a�4�
�;�}�W���*����|!��d��Uʥ�b��<�&�2�h�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����lQ��V��*���
�%�#�1�m��W���&����p]ǻN��*݊�4�;�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����t��D1��C���
�9�u�u���3���>����F�G1��2���&�0�b�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�N����]��hY�����1�o��u���8���B�����h)�����
�u�u����;���:����g)��]����!�u�|�_�w�}�(؁�����V9��V�����u������4�ԜY�Ƽ�9��^ ����o��u����>���<����N��
�����e�n�u�u�'�j�0���
����l��A��Oʜ�u��
���f�W���	�ߓ�Z��[��*���u������4�ԜY�Ƽ�
9��P �����e�4�
�9�w�}�9ύ�=����z%��N������2�4�&�2�l�Mϗ�Y����)��tUךU���
�
�<�;�;��(ށ�	����\��yN��1�����_�u�w��(�������V9��N��U���
���n�w�}����*����_��h\�����1�o��u���8���B�����1�����;�&�0�e�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	����`��X�����e�4�
�9�w�}�9ύ�=����z%��N����
�0�%�<�#��(���Y����g"��x)��*�����}�d�3�*����P���F��^�����<�!�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�d��-����&����z(��c*��:���
�����l��������l�N��Dۊ�;� �&�0�g�<�(���Y�ƅ�5��h"��<��u�u�%�d��3�������/��d:��9�������w�n�W������]ǻN��*����%�!�
����������}F��s1��2���_�u�u�
�f�����&����	F��=��*����
����u�FϺ�����O��N����
�;� �&�2�o��������z(��c*��:���n�u�u�%�f�����
����\��yN��1��������}�D�������V�=N��U���d��%�!���(������/��d:��9����_�u�u��l�>�������F��~ ��!�����
����_������\F��d��Uʥ�d�
�;� �$�8�C���&����	F��=��*����n�u�u�'�l�(�������lS�'��&���������W��Y����G	�UךU���
�d��%�#��(ځ�	����\��yN��1�����_�u�w��F���	����V9��N��U���
���
��	�%���Hӂ��]��G�U���%�d�
�;�"�.��������WF��~ ��!�����u�n�2�9�}�������V��E�����u�3�8�g�g�n�1���Y���F�V�����0���
���6���7����|F��d:��;��u�u�4�!�>�(�ϝ�+����}#��c'��*����:�u�0�6�}�W�������G����U���w�e��c�c�;�Gö�
����V��hZ��=��������`����5����c3��q"��!��������/���I߮��l/��b:��4���-�b�e�e�;�i�C��1����}6��h-��6��`�e�e�e�{��(���,����p.��C��Ɲ�������E���L����.��h=��*���h�a�y����(���D����.��h=��*���h�y��
���$��A߮��l5��h(��M���y��
����J��L˛�9F������!�4�
�:�$�����&����`2��{!��6��u�d�n�u�w�>�����ƭ�l��D�����
�u�u����>���D����l�N�����;�u�%���)�(���&����`2��{!��6�����u�g�w�2����I����D��^�E��e�e�e�e�g�m�G��I����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�g�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�g�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���g�u�:�;�8�m�W��[����V��^�E��e�e�e�e�f�m�U�ԜY�Ư�]��Y�����
�!�
�&��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�d�e�e�u�W�W�������]��G1��*���
�&�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�w�]�}�W���
������d:��Ҋ�&�
�u�u���8���&����|4�Y�����:�e�u�h�u�m�G��I����V��^�D��e�e�w�_�w�}��������C9��h��*���
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��_�E��e�w�_�u�w�2����Ӈ��`2��C_�����l�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��_�����e�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��\�����d�o�����4���:����T��S�����|�o�u�e�g�m�G��I����W��^�E��e�n�u�u�4�3����Y����g9��]�����g�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��Z�����f�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��[�����a�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��X�����`�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��Y�����c�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��V�����b�o�����4���:����T��S�����|�o�u�e�g�m�G��H����V��^�E��e�n�u�u�4�3����Y����g9��W�����m�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��^�����l�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��_�����e�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��\�����d�o�����4���:����T��S�����|�o�u�e�g�m�F��I����V��^�E��e�n�u�u�4�3����Y����g9��]�����g�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��Z�����f�o�����4���:����T��S�����|�o�u�e�g�l�G��I����V��^�E��e�n�u�u�4�3����Y����g9��[�����a�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��X�����`�o�����4���:����T��S�����|�o�u�e�f�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��Y�����c�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��V�����b�o�����4���:����T��S�����|�o�u�d�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����\��h��G��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D��ۊ�u�u��
���(���-���F��@ ��U���o�u�d�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�e�l�}�WϽ�����GF��h�����#�g�f�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�f�f�W�������R��V�����
�#�g�c�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�f�m�L���YӅ��@��CN��*���&�
�#�g��g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�F��Y����\��V �����:�&�
�#�e�j�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�F��B�����D��ʴ�
�:�&�
�!�o�O��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�E���Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��H���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��Y��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�D���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�d�w�_�w�}��������C9��Y����
�f�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�e�d�l�}�WϽ�����GF��h�����#�g�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�g��}���Y����G�������!�9�f�
��g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�m�F��Y����\��V �����:�&�
�#�e�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�C��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�E���Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����W��UךU���:�&�4�!�6�����&����lU��-��C��������4���Y����W	��C��\��u�e�d�d�f�m�G��H����W��^�D��e�n�u�u�4�3����Y����\��h��G���`��e�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��H����W��_�D��e�e�e�e�g��}���Y����G�������!�9�f�
���6���Cӵ��l*��~-��0����}�d�1� �)�W���C���W��_�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����A���5��h"��<������}�w�2����I����D��^�E���_�u�u�:�$�<�Ͽ�&����G9��]��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������V��T��!�����
����_������\F��T��W��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�d��i�G��*����|!��h8��!���}�a�1�"�#�}�^��Y����W��^�E��w�_�u�u�8�.��������]��[��3���u��
����2���+����W	��C��\��u�d�d�d�f��}���Y����G�������!�9�d�
�g�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��u�u�6�;�#�3�W�������l
��1�E��������4���Y����W	��C��\��u�e�e�e�f�m�G��I��ƹF��X �����4�
�:�&��+�B��I����g"��x)��*�����}�a�3�*����P���V��_�E��e�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��S�����|�o�u�e�g�m�G��[���F��Y�����%�6�;�!�;�l�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�e�w�_�w�}��������C9��Y����
��o����0���/����aF� N�����u�|�o�u�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��q(��Oʆ�������8���H�ƨ�D��^��O���d�d�d�d�f�l�F��H����F�T�����u�%�6�;�#�1�D݁�I����V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����9��N��1��������}�FϺ�����O�
N��E��u�u�6�;�#�3�W�������l
��h_��U���
���
��	�%���Y����G	�N�U��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�d�w�_�w�}��������C9��Y����
�g�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�e�e�l�W�W���������t=�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E���_�u�u�!�%�?����
����P	��Y	��U���<�2�_�u�w�)�����ƪ�^9��T�����3�4�
��1�0�Mϭ�����Z�Y��W�ߊu�u�<�;�;�<�(���&����l5��D�����e�o�����4�ԜY�ƿ�T�������7�1�a�u�w��;���B�����Y������;�4��9�/����I����@��N��1�����_�u�w�4����	�ғ�R��[-�����
�
�
�'�0�g�$���5����\�^�����u�<�;�9�'�i�:�������G��h��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�a��9�<�4�������lV��G1�����0�u�u����>���D����l�N�����u�
�
�4�"�1��������9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������]��[1��D���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W�������lR��V �����!�:�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�M����F��X �����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����R
��Y�����g�<�
�<�w�}�#���6����9F������%�a��;�6���������l��PN�&������o�w�m�L���Yӕ��]��G1��8���4��;�'�;�8�E���&����Z��^	��U���
���n�w�}�����Ƽ�9��Y��6���'�9�0�g�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l+��B�����:�
�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*��� �9�:�!�8��(܁����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�a��3��������l��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�a��;�4��3�����Փ�C9��S1�����u��
���}�J���^���F��P ��U���
�4� �9�8�)����&ǹ��l��T��!�����n�u�w�.����Y����~��V�����9�0�a�%�2�}�W���&����pF��I�N���u�&�2�4�w��(�������]��[1��A���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�6�(��������V9��V�����'�2�o����0���C���]ǻN�����9�%�a��9�<�4�������lS��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������\��X��*ߊ�'�2�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�l�}�Wϭ�����C9��z�����;�'�9�0�b�<�(���&����Z�=��*����n�u�u�$�:����&ǹ��]��t�����0�`�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�M����F��X �����
�
�;�&�0�g�$���5����l�N�����u�
�
�4�"�1��������9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*��� �9�:�!�8��(ف�	����l��D��Oʆ�����]�}�W�������lR��V �����!�:�
�
��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��Y��6���'�9�0�b�>�����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��A���;�4��;�%�1����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
��<��������_9�� 1��*���
�;�&�2�m��3���>����F�D�����
�
�4� �;�2����&����R��[
�����o������M���I��ƹF��^	��ʥ�`��;�0�2�m��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�`��;�0�2�m����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�
�
�4�0��(߁�	����l��D��Oʆ�����]�}�W�������lS��V ��*���
�%�#�1�'�8�W���-����t/��S��E��u�u�&�2�6�}�(ځ�����V9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(ځ�����V9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�>�3�Ϯ�L����T��h_�����1�<�
�<�w�}�#���6����9F������%�`��;�2�8�F���&����C��T��!�����u�h�p�z�}���Y����R
��h[�����
�
�
�;�$�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h[�����
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��@���;�0�0�g�6���������\��c*��:���n�u�u�&�0�<�W���&����V9��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�`��3����J����@��N��1��������}�D�������V�=N��U���;�9�%�`��3����J����TF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���&�2�4�u������&����R��[
�����2�o�����4�ԜY�ƿ�T����*���2�
�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����a��R1��A���
�<�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����a��R1��A���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W�������lS��V ��*���
�%�#�1�>�����Y����)��tUךU���<�;�9�%�b������ғ�C9��S1�����u��
���}�J���^���F��P ��U���
�4�2�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�4�2�
������Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������%�`��;�2�8�B���&����Z��^	��U���
���n�w�}�����Ƽ�9��Y	�����4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�B�������lP��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�B�������lP��E��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�&�0�<�W���&����V9��1��*���
�;�&�2�m��3���>����F�D�����
�
�4�2���(�������A��N��1�����o�u�g�f�W���
����_F��1�����0�b�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����0�b�%�0�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�ƿ�T����*���2�
�
�
�'�+����&����	F��s1��2���_�u�u�<�9�1����+����l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
�6�:�(���&����Z�=��*����
����u�FϺ�����O��N�����4�u�
�
�6�:�(���&����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���<�;�9�%�b������ޓ�C9��S1��*���u�u��
���L���Yӕ��]��G1��'���0�0�m�4��1�(�������g"��x)��U��r�r�_�u�w�4����	�ӓ�R��h��*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�ӓ�R��h��*���2�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�n�w�}�����Ƽ�9��Y	�����4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
��<����&ʹ��l��h���������g�W��B�����Y������'�8�!�%��(߁�����\��c*��:���
�����l��������l�N�����u�
�
�4�6�8�����֓�A��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�&�2�4�w��(�������A��h^�����1�<�
�<�w�}�#���6����9F������%�c��'�:�)����&ù��l��h���������g�W��B�����Y������'�8�!�%��(ށ�����\��c*��:���
�����l��������l�N�����u�
�
�4�6�8�����ד�A��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�&�2�4�w��(�������A��h_�����1�<�
�<�w�}�#���6����9F������%�c��'�:�)����&¹��l��h���������g�W��B�����Y������'�8�!�%��(܁�����\��c*��:���
�����l��������l�N�����u�
�
�4�6�8�����Փ�A��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�&�2�4�w��(�������A��h]�����1�<�
�<�w�}�#���6����9F������%�c��'�:�)����&����l��h���������g�W��B�����Y������<�&�0�g�4�(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������<�&�0�g�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����
�
�4�;���(�������]9��PN�&������_�w�}����Ӗ��l!��Y��*ڊ�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��(�������9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1����>����l��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�b��<�&�2�l��������V�=��*����u�h�r�p�W�W���������h)�����
�
�;�&�0�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h)�����
�
�'�2�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�L���Yӕ��]��G1��2���&�0�g�4��1�(���
���5��h"��<��u�u�&�2�6�}�(؁�����V9��V�����'�2�o����0���C���]ǻN�����9�%�b��>�.��������TF��d:��9�������w�n�W������]ǻN�����9�%�b��>�.����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
��<����&����l��h�����o������}���Y����R
��hY�����
�
�
�%�!�9����Y�Ɵ�w9��p'��O���e�n�u�u�$�:����&Ĺ��Z��R1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&Ĺ��Z��R1�����u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}����Ӗ��l!��Y��*ފ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�b��4����M����E
��G��U����
���w�`�P���s���@��V��*݊�4�;�
�
��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*݊�4�;�
�
��/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʥ�b��<�&�2�h��������l��T��!�����n�u�w�.����Y����t��D1��@���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�j�0���
����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�j�0���
����l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�&�2�6�}�(؁�����V9��V�����;�&�2�o���;���:���F��P ��U���
�4�;�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��p�����b�<�
�<�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��p�����b�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����R
��hY�����
�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�@�������lQ��G1�����0�u�u����>���D����l�N�����u�
�
�4�9��(ׁ�����\��c*��:���
�����l��������l�N�����u�
�
�4�9��(ׁ����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�b��4����A����E
��^ �����u��
���f�W���
����_F�� 1�����0�m�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�N����]��hW�����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�N����]��hW�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����t��D1��L���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�6�3�(���&����_��E��Oʆ�����m�}�G��Y����Z��[N��L���2�4�&�0�g�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�d�$�������lV��E��Oʆ�����m�}�G��Y����Z��[N��L���2�4�&�0�g�<�(���&����Z�=��*����n�u�u�$�:����&ʹ��T��D1��E���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�d�$�������lW��Y1���������W�W���������h=�����
�
�
�'�0�g�$���5����\�^�����u�<�;�9�'�d�$�������lW��G1�����
�<�u�u���8���B�����Y������2�4�&�2�l��������V�=��*����u�h�r�p�W�W���������h=�����
�
�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�>�3����&����V�=��*����u�h�r�p�W�W���������h=�����
�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�N�������l��h�����%�0�u�u���8���Y���A��N�����4�u�
�e��)����
����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�l�(���	����@9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	����`��X�����e�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u��m�$�������l��h�����%�0�u�u���8���Y���A��N�����4�u�
�d��-����&ù��l��T��!�����
����_������\F��d��Uʦ�2�4�u�
�f�����&����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�<�;�;�-�Fށ�����l��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�d�
�;� �$�8�G���&����C��T��!�����u�h�p�z�}���Y����R
��h_��<���!�
�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����D���%�!�
�
��/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʥ�d�
�;� �$�8�F���&����Z��^	��U���
���n�w�}�����Ƽ�W��Y�����d�4�
�9��/���*����|!��T��R��_�u�u�<�9�1���&����G��h\�����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�H¹��C��h��*���2�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�n�w�}�����Ƽ�W��Y�����g�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u��l�>�������9��h��*���2�o�����4��Y���9F������%�d�
�;�"�.��������TF��d:��9�������w�n�W������]ǻN�����9�%�d�
�9�(����J����TF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���&�2�4�u��l�>������� 9��h��*���&�2�o����0���s���@��V��*����%�!�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��h'�� ���0�a�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��_�����&�0�a�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*����%�!�
����������@��N��1�����_�u�w�4����	����z��C��*ފ�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��F���	����V9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(���0����@9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	����z��C��*ߊ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�d��3�����ӓ�C9��S1�����u��
���}�J���^���F��P ��U���d��%�!���(���
���5��h"��<������}�f�9� ���Y����F�D�����
�d��%�#��(ف����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�d��3�����Г�C9��S1��*���u�u��
���L���Yӕ��]��G1�*��� �&�0�c�6��������5��h"��<���h�r�r�_�w�}����Ӆ��u#��u/����� �
�l�e�2�m�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����Y�����3�
�g�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hY�U����
�����#���Q����\��XN�N���u�&�2�4�w�-��������`2��CZ�����u�u��
���L���Yӕ��]��V�����1�
�d�u�w��;���B�����Y�����<�
�&�$���؁�
����	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��R��!���d�
�&�
�f�g�$���5����l�N�����u�%�&�2�5�9�B��CӤ��#��d��Uʦ�2�4�u�'��(�@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʧ�2�b�d�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l �� Z�����u��
����2���+������Y��E��u�u�&�2�6�}����A����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��Z�Oʗ����_�w�}����Ӂ��l ��h��D���
�d�
�%�3�3�W���-����t/��=N��U���;�9�4�
�>�����*����
9��Z1�Oʆ�����]�}�W�������C9��P1�����`�o�����}���Y����R
��G1�����0�
��&�f�����J����g"��x)��N���u�&�2�4�w�-��������R�,��9���n�u�u�&�0�<�W���&����U9��h��C���4�
�:�0�m��3���>����F�D�����
�
�<�;�;��(݁�����V��Q��L؊�g�o�����4���:����V��X����n�u�u�&�0�<�W���
����@��d:�����3�8�g�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��e�W���6����}]ǻN�����9�4�
�<��.����&����l ��h\�Oʆ�����]�}�W�������C9��P1�����e�o�����}���Y����R
��E�� ��m�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����_��N��1��������}�D�������V�=N��U���;�9�2�%�1��B܁�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�e�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U��Y��G��������4���Y����W	��C��\�ߊu�u�<�;�;�/���@����g"��x)��*�����}�d�3�*����P���F��P ��U���
�d�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z��D��&���!�b�3�8�f�}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(�������@��h��*��o������}���Y����R
��G1�����1�c�c�o���2���s���@��V�����2�7�1�b�`�g�5���<����F�D������-� ��9�(�(���H����V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�1��:���K����lT��1����e�u�u����>���<����N��
�����e�n�u�u�$�:����*����2��x��Gڊ�
� �d�l��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1�� ���;� �
�e�d�/���I����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʶ�
�����(����Lʹ��9��P1�D���u��
����2���+������Y��E��u�u�&�2�6�}��������l��N��1��������}�D�������V�=N��U���;�9�3�
���8���H¹��A��Y�U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���N�ѓ�F��d:��9�������w�n�W������]ǻN�����9�3�
������&¹��T9��]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��3��������Z��D=�����e�'�2�d�e�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h �����'�
�<�6�$�����H����lW��N�&���������W��Y����G	�UךU���<�;�9�3���;�������_��[��B���3�
�c�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��O#��!���!��9�<�;��@�������R��N��1��������}�D�������V�=N��U���;�9�3�
������&����Z��h_��D���
�c�
�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��b"��:����9�<�9��i�F�������F��d:��9�������w�n�W������]ǻN�����9�3�
���$��������_��h_�����b�g�o����0���/����aF�N�����u�|�_�u�w�4��������T9��R��!���d�
�&�
�w�}�#���6����9F������4�
�<�
�3��F���Y����v'��=N��U���;�9�3�
������&����Z��h_��D���2�d�`�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l��{:�� ��� �!�%�,�a�l����H����	F��s1��2������u�d�}�������9F������3�
���.�(�(�������lW��1����c�u�u����>���<����N��
�����e�n�u�u�$�:����*����w��C1�*ۊ�0�
�b�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�d�
�$��E��*����|!��d��Uʦ�2�4�u�%�$�:����A���$��{+��N���u�&�2�4�w����� ����`��E��*���d�'�2�d�`�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h �����'�
�=�0��<����&����9��P1�M���u��
����2���+������Y��E��u�u�&�2�6�}��������A��_��%���0��
�'������N���5��h"��<������}�f�9� ���Y����F�D������;�1�
�2�0�#�������V6��h��*���
�b�c�o���;���:����g)��]����!�u�|�_�w�}����Ӆ��]	��h�����&�4�0��9�/��������V��N��1��������}�D�������V�=N��U���;�9�4�
�>�����*����S��D��A�������W�W���������D�����m�d�o����9�ԜY�ƿ�T��	��*���
�
�
� �a�i�������5��h"��<��u�u�&�2�6�}��������A��V�����:�!�:�
������A���5��h"��<������}�f�9� ���Y����F�D�����9�;�1�
�2�0�4�������\��X��*؊�0�
�m�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������_9��S������&�4�0��3����
�Փ�V��_�Oʆ�������8���J�ƨ�D��^����u�<�;�9�4���������p��V
��6���'�9�&�a�%�:�F��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����:�0�!�'��<��������A	��D1�����d�g�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����\��C��*���6�1�1�:�#�2�(���&����^��T��!�����
����_������\F��d��Uʦ�2�4�u�9�9�9�(�������P��S-�����
�
�
�0��e�@��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������
�0�8��$�<��������l��h��*��g�o�����4���:����U��S�����|�_�u�u�>�3�Ͻ�&����l��Z1�����0��;�'�;�.�N�������F��d:��9�������w�n�W������]ǻN�����9�3�
���	����I�ԓ�F9�� W��F��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���<����G9��h\�����m�a�o����0���/����aF�N�����u�|�_�u�w�4��������#��x��B܊�
� �d�m��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1��9����!�b�
��8�(��I����g"��x)��*�����}�d�3�*����P���F��P ��U���&�2�6�0��	���&����_�=��*����n�u�u�$�:����	����l��hV�U������n�w�}�����ƪ�l��u�����'�2�d�c�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��z;��G���!�b�d�3��i�E���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�������g��#�j�F�������F��d:��9�������w�n�W������]ǻN�����9�3�
��/�(�(�������_��N�&���������W��Y����G	�UךU���<�;�9�4��4�(�������@��h��*���o������}���Y����R
��G1�����1�m�m�o���2���s���@��V�����
�
�
�
�"�k�C���&����GF��d:��9����_�u�u�>�3�Ϲ�	����l ��h��C���4�
�1�0�m��3���>����F�D�����'�
�
�
�����M����A��NN�&������_�w�}����Ӂ��l ��h��*���c�a�<�
�6�:�(؁�&����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�e�3�d�;�(��&����R��hY��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù�� 9��hX�*����;�0�b�2�o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �c�c�4�(�������V9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������9��h<�����
�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����a�
�;��9�8�@���L����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�A�������]�� 1��C��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����l ��Z�����4�2�
�
��}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���f�3�
�a��3�:�������G��h_����o������}���Y����R
��E��*ڊ�
�
� �c�c�4�(�������]��[1�*���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����U9��Q��Aފ�;��;�4��3����H����F��d:��9����_�u�u�>�3�Ϲ�	����l ��h��C���<�
�4� �;�2����&�ԓ�lU�=��*����
����u�FϺ�����O��N�����4�u�'�
���(܁�����l��z�����;�'�9�d���W���-����t/��=N��U���;�9�2�%�1�m��������9��h#�� ���:�!�:�
�e�8�B��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���
�
�
� �a�i��������p	��E��D؊�
�u�u����>��Y����Z��[N�����e�3�f�3��i�(���4����_%��C��*���0�b�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h]�� ��a�<�
�4�9��(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�e�3�f�1��Cہ�����]��h��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����U��Z�����<�&�a�0�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���
� �c�a�>�����&ǹ�� F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�D���&����Z��V��*ފ�
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�;��<�$�i���Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
�
�
�"�k�C���&����@9��R1�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-�����Փ�F9��1��*���;�
�
�
�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q1�����3�
�a�
�9�/����I����g"��x)��N���u�&�2�4�w�/�(���&����U��Z�����
�
�
�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��1��F���
�a�
�;���(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�e�3�f�1��Cہ�����9��N�&���������W��Y����G	�UךU���<�;�9�2�'�;�G���J����R��^ ��#���0�f�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h]�� ��a�<�
��f�8�G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���
�
�
� �a�i����)�ד�lW�=��*����
����u�FϺ�����O��N�����4�u�'�
���(܁�����l��E�����u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����U9��Q��Aފ�%�'�!�'��}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���f�3�
�a��-��������	F��s1��2������u�d�}�������9F������2�%�3�e�1�n����Mǹ��l��B��F��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����l ��Z�����0� �;�a�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��h^��*ي� �c�a�4��8����L����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�A�������G��hX��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��(߁�&����lP��h�����'�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����a�
�%�'�#�/�(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�f�3��i�(�������]9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������9��h��Oʆ�����]�}�W�������A��h^��*���3�
�l�
�'�.����Cӵ��l*��~-�U���&�2�4�u�%��(߁�&�ԓ�F9��1��*���0�o�����4�ԜY�ƿ�T��	��*���
�
�g�3��d�(�������\��c*��:���n�u�u�&�0�<�W���&����U9��h��C���<�
��'�9�8�N���I����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
�e�;�(��&����*��Y	��L���d�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����l ��1��*��
�;�'�&�#�i�Mύ�=����z%��N�����4�u�'�
���(�������
9��h>�����&�m�0�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��h^��*���3�
�l�
�9��;�������V9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m���&����
_��Y1�����;�e�0�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��h^��*���3�
�l�
�9�����	����W ��F1�U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����l ��W������`�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h_�����l�
�;���}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���d�
� �c�n�<�(�������\��c*��:���
�����l��������l�N�����u�'�
�
���E���&����R��R����o������!���6���F��@ ��U���_�u�u�<�9�1�����֓�lW��Q��Lӊ�%�'�!�'��}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���d�
� �c�n�<�(�������\��c*��:���
�����l��������l�N�����u�'�
�
���E���&����R��RN�&������_�w�}����Ӂ��l ��h��D���
�d�
�%�$�<���*����|!��d��Uʦ�2�4�u�'���(���H����W��V�����o������}���Y����R
��E��*ڊ�
�d�3�
�f��������5��h"��<��u�u�&�2�6�}����&ù��W��B1�C���
�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�*���b�c�4�
�2�(���Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
�
�d�1��Fف�	����F��N�&���������W��Y����G	�UךU���<�;�9�2�'�;�G���H¹��lQ��h�����u��
���f�W���
����_F��G1��E���f�3�
�a��-��������@��C1���������g�W��B�����Y�����3�e�3�d��(�A�������R��V�����
�0�u�u���8���Y���A��N�����4�u�'�
���(�������9��h�����%�&�4�!�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�<�(���&����l5��D�*���
�b�o����0���s���@��V�����2�7�1�d�b�}�W���5����9F������2�%�3�
�e��G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���b�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�l��h�����
�!�
�&��}�W���&����p]ǻN�����9�4�
�<��9�(��L����|)��v �U���&�2�4�u�'�.��������l��h��*���u��
���f�W���
����_F��h��*���
�e�g�o���2���s���@��V�����2�6�0�
��.�Fށ�
����\��c*��:���n�u�u�&�0�<�W���
����W��Y�Oʗ����_�w�}����Ӈ��@��T��*���&�d�
�&��j�Mύ�=����z%��N�����4�u�%�&�0�?���A����q)��r/�����u�<�;�9�6�����
����g9��\�����d�o�����4�ԜY�ƿ�T�������7�1�d�l�w�}�8���8��ƹF��^	��ʲ�%�3�
�g��m�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U��]��E��������4���Y����W	��C��\�ߊu�u�<�;�;�:����&����CW�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�j�@���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�
�f�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��B���%�u�u����>���<����N��
�����e�n�u�u�$�:��������lQ��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-����M˹��\��c*��:���
�����l��������l�N�����u�'�
� �`�e����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�`�
�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��B1�F���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����Q��N�&���������W��Y����G	�UךU���<�;�9�2�'�;�(��&���5��h"��<������}�f�9� ���Y����F�D������-� ���)�:�������Q��h��B���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����2��B�� ���%�,�d�
��(�@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
���,�"�����	����9��Q��C܊�e�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����g��C1�����9�
�a�d�1��Aف�H����g"��x)��*�����}�d�3�*����P���F��P ��U���4�g�&�3��o�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
� �m�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������
��h8��L���
�f�
�d�m��3���>����v%��eN��Gʱ�"�!�u�|�]�}�W�������^��h��*���3�
�a�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��^1�����
�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƾ�G9��^1�����`�
�f�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lW��h��*��� �m�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�����
�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G\��*���m�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӕ��lT��h��*���!�6�&�
�"�e�B���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����!�%�<�3��j�(��Cӵ��l*��~-��0����}�a�1� �)�W���s���@��V��*��� �!�m�
�"�d�F���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�������g��#�o�(�������lW��B1�L���u�u��
���(���-���Q��X����n�u�u�&�0�<�W���&����l_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��G߁�&����W��N�&���������W������\F��d��Uʦ�2�4�u�8��(�N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�f�3�
�c��D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��D���3�
�a�
�f�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��_�� ��f�%�u�u���8���&����|4� N�����u�|�_�u�w�4����	����9��^1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������9��Q��Cۊ�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�+����G9��h��L���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����2��x��Gڊ�;�3��%��(�O���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʦ�9�!�%�
��(�N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�b�<�1��Nށ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�
�"�d�@���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��&��� ��;� ��m����A¹��\��c*��:���
�����l��������l�N�����u�
�4�g�`����H¹��\��c*��:���
�����l��������l�N�����u�:�
�
�g�;�(��L����	F��s1��2������u�`�9� ���Y����F�D�����:�
�
�d�1��G���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʡ�%�<�<�<��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�<�<�<��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʧ�!�<�<�<��(�F��&���5��h"��<������}�c�9� ���Y����F�D�����8�
�f�
���O���&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�ہ�����9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(�������Q��N�&���������W������\F��d��Uʦ�2�4�u�0���(���@����G9��D�� ��`�
�f�o���;���:����g)��_����!�u�|�_�w�}����ӕ��l��h�����e�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�a��[��L���
�e�d�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����U5��z;��G���!�g�
�;�2�-�!�������
_��N�&���������W��Y����G	�UךU���<�;�9�!�'�4�(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�d�g�4�(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�m��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�c�
� �f�n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����m�3�
�d�n�-�W���-����t/��a+��:���b�1�"�!�w�t�}���Y����R
��Z��F���
�d�f�%�w�}�#���6����e#��x<��Bʱ�"�!�u�|�]�}�W�������lV��1��ۊ� �d�g�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hY��ۊ� �d�`�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������R����
� �d�`��h�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1�� ���;� �
�e�>������ד�F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	Ź��l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}�����ѓ�9��h_�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������ZW��B1�M݊�g�o�����4���:����V��X����n�u�u�&�0�<�W���������C1�*؊� �d�b�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��d+��6���!�m�
�
�"�l�@ց�I����g"��x)��*�����}�u�8�3���B�����Y�������� ��k�E���&����l��N��1��������}�GϺ�����O��N�����4�u�
�4�e�e�(���H����CW�=��*����
����u�FϺ�����O��N�����4�u�:�
��o����K�ғ�F��d:��9�������w�j��������l�N�����u�:�
�
�d�;�(��M����	F��s1��2������u�e�}�������9F������!�%�<�<�>��N���&����l��N��1��������}�GϺ�����O��N�����4�u�8�
���F���&����l��N��1��������}�GϺ�����O��N�����4�u�0�
���F���&����l��N��1��������}�F�������V�=N��U���;�9�!�%�f�l����¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&�ӓ�F9��^��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���K����U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�/��������W��V�����
� �d�f��n�Mύ�=����z%��r-��'���a�1�"�!�w�t�}���Y����R
��R�����`�3�
�f�e�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1�����
�
� �d�`��D��*����|!��h8��!���}�b�1�"�#�}�^�ԜY�ƿ�T��������;� �
��3����/�ד�F9�� V��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)����&���� ^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�l�@�������
V��N�&���������W������\F��d��Uʦ�2�4�u�8��i����J�Г�F��d:��9�������w�m��������l�N�����u�8�
�`�1��C���	����`2��{!��6�����u�b�3�*����P���F��P ��U���
�d�
� �f�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �d�g��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��\�*ۊ�g�3�
�a�e�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��C��M݊�
� �d�f��n�Mύ�=����z%��r-��'���e�1�"�!�w�t�}���Y����R
��h<�� ���l�
� �d�d��B��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��������;� �
��3����	����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�(���O����U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	Ĺ��l ��Z�*��o������!���6�����Y��E��u�u�&�2�6�}�����ޓ�9��h_�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����4����])��hY�� ��`�
�d�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��}#��x��Dڊ�:�<�!�<�1��C���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
��-� ��m��������R��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-����Kƹ��P	��T��!�����
����_�������V�=N��U���;�9�2�%�1��Eځ�����g"��x)��N���u�&�2�4�w�-��������`2��CX�����u�u��
���L���Yӕ��]��V�����1�
�`�g�m��8���7���F��P ��U���&�2�6�0��	���&����S�=��*����n�u�u�$�:����	����l��h_�D������]�}�W�������C9��P1������&�d�
�$��O��*����|!��d��Uʦ�2�4�u�%�$�:����H����	F��x"��;�ߊu�u�<�;�;�:����&����\��S��U���
���
��	�%���Y����G	�UךU���<�;�9�2�'�;�(��&���5��h"��<��u�u�&�2�6�}��������l��N��1�����_�u�w�4��������F9�� 1��U����
���l�}�Wϭ�����R��d1����������4���Y����W	��C��\�ߊu�u�<�;�;�<�(���&����T��N��:����_�u�u�>�3�Ͽ�&����Q��Z�Oʗ����_�w�}����Ӈ��@��U
��A��o�����W�W���������D�����a�`�o����9�ԜY�ƿ�T�������7�1�a�a�m��8���7���F��P ��U���&�2�7�1�c�n�MϜ�6����l�N�����u�%�&�2�5�9�C��CӤ��#��d��Uʦ�2�4�u�%�$�:����L���$��{+��N���u�&�2�4�w�-��������R�,��9���n�u�u�&�0�<�W���
����W��]��U�����n�u�w�.����Y����Z��S
��G���u����l�}�Wϭ�����R��^	�����f�u�u����L���Yӕ��]��V�����1�
�a�u�w��;���B�����Y�����<�
�1�
�c�}�W���5����9F������4�
�<�
�3��B���Y����v'��=N��U���;�9�4�
�>�����O����q)��r/�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��S1�A������]�}�W�������C9��P1����f�o�����}���Y����R
��G1�����1�g�g�o���2���s���@��V�����2�7�1�g�f�g�5���<����F�D�����%�&�2�7�3�o�G��;����r(��N�����4�u�%�&�0�?���@����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lT��T��:����n�u�u�$�:����	����l��h\�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�l�u�u���6��Y����Z��[N��*���
�1�
�d�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&���� R��N��:����_�u�u�>�3�Ͽ�&����Q��[�Oʗ����_�w�}����Ӈ��@��U
��F��o�����W�W���������D�����f�`�o����9�ԜY�ƿ�T�������7�1�f�a�m��8���7���F��P ��U���&�2�7�1�d�n�MϜ�6����l�N�����u�%�&�2�5�9�C��CӤ��#��d��Uʦ�2�4�u�%�$�:����M���$��{+��N���u�&�2�4�w�-��������V�,��9���n�_�u�u�8�-����Y����P��q��*���u��u�u�'�/�W�ԜY���F��h��U���������}���Y���R��D��U��������W�W���Y�ƭ�l��E��U��������W�W���Y�ƭ�l��RN�:��������W�W���Y�ƭ�l��RN�:��������W�W���Y�ƭ�l��S��U���u��
���f�W���Y����]9��Y	��B���e�o��u���8���&����|4�_�����:�e�n�u�w�}�WϷ�&����V9��R1�Oʜ�u��
����2���+������Y��E��u�u�u�u�>�����&Ĺ��F��~ ��!�����
����_������\F��d��U���u�<�
�4�0��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����4�2�
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h<�����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����R��hY��*���u������4���:����U��S�����|�_�u�u�w�}��������l��T��;ʆ�������8���J�ƨ�D��^����u�u�u�;��3��������lW��R1�Oʜ�u��
���f�W���Y����]9��Y��6���'�9�d�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h#�� ���:�!�:�
�e�8�E��0�Ɵ�w9��p'�����u�u�u�;��3��������lW��R1�Oʜ�u��
����2���+������Y��E��u�u�u�u�>���������A	��\��*���u������4�ԜY���F��h#�� ���:�!�:�
�e�8�B��0�Ɵ�w9��p'��#����u�f�u�8�3���B���F���8���4��;�'�;�l�(���Y�ƅ�5��h"��<��u�u�u�u�>���������A	��\��*���u������4���:����U��S�����|�_�u�u�w�}��������l��T��;ʆ�������8���J�ƨ�D��^����u�u�u�;��4�������/��d:��9�������w�n�W������]ǻN��U���;��<�&�c�8�E��0�Ɵ�w9��p'��#����u�f�u�8�3���B���F���2���&�a�0�f�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����]9��^ ��A���a�o��u���8���&����|4�_�����:�e�n�u�w�}�WϷ�&����@9��R1�Oʜ�u��
����2���+������Y��E��u�u�u�u�>�����&ǹ��F��~ ��!�����
����_������\F��d��U���u�<�
�4�9��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����0�0�
�u�w��$���5����l�N��Uʼ�
��g�0�g�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Y�����g8��*���u�u�����0���/����aF�N�����u�|�_�u�w�}�W���)����V9��N��U���
���
��	�%���Hӂ��]��G�U���u�u�<�
��o���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N�����
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƥ�l5��1��D���u��
���(���-��� W��X����n�u�u�u�w�<�(�������\��b:��!�����
����_������\F��d��U���u�4�
�0�"�3�F��6����g"��x)��*�����}�d�3�*����P���F�N��*��� �;�g�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƭ�l��B��F��������4���:����U��S�����|�_�u�u�w�}��������F��x;��&���������W��Y����G	�UךU���u�u�%�'�#�/�(���Y����`2��{!��6�����u�f�w�2����I��ƹF�N�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����C9��C��*���u� �u����>���<����N��
�����e�n�u�u�w�}��������l^�!��U���
���
��	�%���Hӂ��]��G�U���u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�N�����0�o��u���8���Y��ƹF��Y
�����;�;�n�_�w�}����������s^�A���e�3�d�u��}�WϮ����F�N�����9�u�u����;���:���F�N��*���u�u�����0���s���F�V�����u�u�����0���s���F�V�����o������0���s���F�V�����o������0���s���F�V�����u�u� �u���8���B���F���%���4�2�
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h>�����0�l�0�d�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����]9��D��A���u��
���L���Y�����g"�����
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƥ�l6��P�����0�d�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������R��Y1����o��u����>���<����N��
�����e�n�u�u�w�}��������C��R
�����`�o��u���8���&����|4�_�����:�e�n�u�w�}�WϷ�&����\��yN��1��������}�D�������V�=N��U���u�;��
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���R��R����o������0���/����aF�N�����u�|�_�u�w�}�W�������]9��N��!ʆ�������8���J�ƨ�D��^����u�u�u�%�%�)����Y�ƃ�gF��s1��2������u�d�}�������9F�N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���Y�����T��U��������t�}���Y����P	��X ���ߠ_�u�u�:�'�3����I���� R��h^��*���_�u�u�8�)�_���Y�����T��Oʜ�u��
���f�W���Y����C9��CN�<����
���l�}�W���YӇ��@��CN�<����
���l�}�W���YӇ��W	��T�� ����
���l�}�W���YӇ��Z��T�� ����
���l�}�W���YӇ��A��NN�:��������W�W���Y�ƥ�l��T��;ʆ�������8���J�ƨ�D��^����u�u�u�%�%�)����Y�ƃ�gF��s1��2������u�d�}�������9F�N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���Y�����T��U��������t�}���Y����P	��X ���ߠ_�u�u�:�'�3����I���� R��h^�����&�7�f�;��o���&����_
��D��&���u�2�;�'�4�u�W���Y����wF��~ ��2���_�u�u�u�w��(���>����z(��p+�����u�u�u�<�g�
�3���Cӯ��v!��d��U���u�1�;�
��	�W���7����a]ǻN��U���:�!����g�>���>���l�N�����_�u�u�u�w�1�W���7ӵ��l*��~-�U���u�u�'�&�#�g�>���-����t/��=N��U���u�<�e�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӂ��F��~ ��!�����
����_������\F��d��U���u�:�6�1�w�}�9ύ�=����z%��r-��'���u�:�;�:�g�f�W���Y����VF��~ ��!�����n�u�w�}�WϺ�����|3��d:��9�������w�n�W������F�=N��U���u�:�%�;�9�f�}���YӅ��C	��Y��Eؑ�c�a�3�e�1�(�(���
����@9��h]�� ���1�%��_�w�}�������F�N��<���u����l�}�W���YӨ��l5��p+��U�����n�u�w�}�WϺ�ù��w2��N��!����_�u�u�w�}����.����\��y:��0��u�u�u�u�3�(�(���-����z(��p+��\�ߊu�u�:�!��}�W���YӅ��\��yN��1�����_�u�w�}�W�������z(��c*��:���n�u�u�u�w�9����Y����g"��x)��*�����}�d�3�*����P���F�N�����u������4���:����U��S�����|�_�u�u�w�}���0�Ɵ�w9��p'�����u�u�u�:�#�g�8���*����|!��h8��!���}�d�1�"�#�}�^���s���V��T�����!�_�_�u�w�2�����ơ�"��Z��*ڊ�8�9�f�;��o���&¹��K9��GN�����u�0�0�<�w�W�W���Y�ƅ�\��y:��0��u�u�u�u���$���<����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�<�d����Mϗ�-����l�N��Uʱ� �
���w�}�9���<���9F������u�u�u�u�3�3�W���7ӵ��l*��~-��0����}�d�1� �)�W���s���F�S��U���������!���6���F��@ ��U���_�u�u�u�w�2���6����g"��x)��*�����}�d�3�*����P����F�R �����:�0�!�_�]�?����Y����A��h^��*ي� �c�a�o�4�0����Ӌ��wV��(��E���f�u�u�%�%�}����s���F�V�����k�4�
�9�{�}�W���YӇ��A��
P�����!�_�u�u�w�}�������F��G1��E���f�3�
�a��-�������F�N��*���0�h�u�'���(���&����R��G1�����u�u�u�u�6�����D�ƫ�C9��1��F���
�a�
�%�>�1�[���Y�����E����u�'�
�
���(���O�ғ�C9��V
�����u�u�u�;��3�������F��G1��E���f�3�
�a��3�%����ѓ�lV�N��U���<�
�4�2���(���GӁ��l ��h��*���c�a�<�
�6�:�(؁�&��ƹF�N�����;�0�b�0�e�`�W���&����U9��Q��Aފ�;��;�0�`�8�E�ԜY���F��h<�����
�
�u�k�0�-�����Փ�F9��1��*���2�
�
�
�{�}�W���Yӏ��a��R1����h�u�'�
���(܁�����l��e�����0�a�_�u�w�}�W���+����lQ��h[��Kʲ�%�3�e�3�d�;�(��&����R��hY��*���u�u�u�u�>�����&Ĺ��F�	��*���
�
�
� �a�i��������9��BךU���u�u�;��9�8�@���N���T��Q1�����3�
�a�
�9�����N����l�N��Uʼ�
�4� �9�8�)����K����[�P�����3�f�3�
�c���������\��X��G���e�_�u�u�w�}��������\��X��G���d�h�u�'���(���&����R��Y1������;�'�9�f��(��Y���F��Y1������;�'�9�f��(���GӁ��l ��h��*���c�a�<�
�6�(��������T��h\�U���u�u�<�
�6�(��������T��h]��Kʲ�%�3�e�3�d�;�(��&����R��[-�����
�g�0�f�]�}�W���Y����R��[-�����
�g�0�a�j�}����&ù�� 9��hX�*����;�4��9�/���&����9F�N��U����;�4��9�/���&����X��E��*ڊ�
�
� �c�c�4�(�������]��[1�*���y�u�u�u�w�4�(�������]��[1�*���u�k�2�%�1�m��������9��h#�� ���:�!�:�
�e�8�A�ԜY���F��h#�� ���:�!�:�
�e�8�@��Y����U9��Q1�����a�
�;��9�<�4�������9�� BךU���u�u�;��>�.�C���I���T��Q1�����3�
�a�
�9�����M����l�N��Uʼ�
�4�;�
���W�������lV��h]�� ��a�<�
�4�9��(���U���F���2���&�a�0�g�j�}����&ù�� 9��hX�*����<�&�a�2�o�}���Y���Z��V��*ފ�
�u�k�2�'�;�G���J����R��^ �����
�
�
�y�w�}�W�������Z��1��A��u�'�
�
���(���O�ғ�]9��^ ��A���a�_�u�u�w�}��������l��S����3�e�3�f�1��Cہ�����]��h��Y���u�u�u�<��<����&����X��E��*ڊ�
�
� �c�c�4�(�������V9��=N��U���u�;��<�$�i���D�ƫ�C9��1��F���
�a�
�;��4��������F�N�����0�0�
�u�i�:����I����l ��Z�����0�0�
�y�w�}�W�������lT��h^��Kʲ�%�3�e�3�d�;�(��&����e9��R1����u�u�u�;���(���Y����A��h^��*ي� �c�a�<���E���H���F�N��*���g�0�g�h�w�/�(���&����U��Z�����
�
�
�y�w�}�W�������lT��h]��Kʲ�%�3�e�3�d�;�(��&����e9��R1����u�u�u�;���(���Y����A��h^��*ي� �c�a�<���F���I���F�N��*���d�0�d�h�w�/�(���&����U��Z�����
�
�
�y�w�}�W�������G��h^��Kʲ�%�3�e�3�d�;�(��&����V��Y1����u�u�u�%�%�)����Y����A��h^��*ي� �c�a�4��8����H���F�N��*��� �;�g�h�w�/�(���&����U��Z�����!�'�
�y�w�}�W�������G��h]��Kʲ�%�3�e�3�d�;�(��&����V��Y1����u�u�u�%�%�)����Y����A��h^��*ي� �c�a�4��8����M���F�N��*��� �;�`�h�w�/�(���&����U��Z�����!�'�
�y�w�}�W�������G��hX��Kʲ�%�3�e�3�d�;�(��&����V��Y1����u�u�u�%�%�)����Y����A��h^��*ي� �c�a�4��8����N���F�N��*��� �;�m�h�w�/�(���&����U��Z�����!�'�
�y�w�}�W�������G��hW��Kʲ�%�3�e�3�d�;�(��&����V��Y1����u�u�u�%�4�}�IϹ�	����l ��h��C���4�
�0�n�]�}�W���&����U9��h��C��o�6�8�:�2�)����I����U9��Q1����u�:�!�8�'�u�W���Y����C9��\N��U���6�>�_�u�w�}�W������F��h��Y���u�u�u�4��)����GӁ��l ��h��G���
�l�
�%�$�<��ԜY���F��h
����u�'�
�
���E���&����R��X �����u�u�u�%�>�1�W�������lV��h_�����l�
�%�<�;�q�W���Y����C9��V
��H���'�
�
�
��o����@ʹ��l��S�U���u�u�<�
��/����@����[�P�����3�d�
� �a�d����5����T��h��Y���u�u�u�<�������ߓ�lW�	N�����e�3�d�
�"�k�N���&����R��hW��*���u�u�u�u�>�����&�����h��*���g�3�
�l��3��������F�N������2�<�&�o�8�G��Y����U9��Q1�*���c�l�<�
��:����A����l�N��Uʼ�
��2�<�$�e���D�ƫ�C9��1��D؊� �c�l�<������
�ޓ�lW�N��U���<�
�!�!���(���Y����A��h^��*���3�
�l�
�9������֓�lV�N��U���<�
�'�1�/�8��������F�	��*���
�
�g�3��d�(���>����K��C�����d�y�u�u�w�}����-���F��G1��E���d�
� �c�n�4�(���L���F�N��*���f�h�u�'���(���K����_��^ ����_�u�u�u�w�-��������X��E��*ڊ�
�g�3�
�n���������JǻN��U���%�'�!�'��}�IϹ�	����l ��1��*��
�%�'�!�%��[���Y�����E�����u�k�2�%�1�m���&����
_��G1�����
�y�u�u�w�}��������lU�	N�����e�3�d�
�"�k�N���&����A��d��U���u�4�
�0�j�}����&ù��T��B1�L���
�0�n�_�w�}����&ù��W��B1�C��6�8�:�0�#�0�E��JǠ��9��_ךU���:�!�8�%��}�W���YӇ��P
��
P�����>�_�u�u�w�}�������R��D�U���u�u�4�
�#�/�W�������lV��h_�����d�
�%�&�6�)�}���Y���R��X ��H���'�
�
�
��l����HŹ��l��RBךU���u�u�%�<�;�}�IϹ�	����l ��1��*��
�%�<�9�{�}�W���YӇ��A��NN��U���
�
�
�
�f�;�(��&����V��d��U���u�<�
�
�w�c�����֓�lW��Q��D܊�;�-�e�_�w�}�W���	����F��N��U���
�
�
�
�f�;�(��&����V��Y1����u�u�u�%�%�)����Y����A��h^��*���3�
�d�
�'�/����&��ƹF�N�����u�k�2�%�1�m���&����P��G1��\�ߠu�u�3�e�1�9����&�Ԣ�lU��D1�*ي� �9�1�%��k�MϽ�����]��\��C���3�e�3�1�1�(�(���
����@9��h]�� ���1�%�u�u�0�3�������9F�N��U���h�u�y�u�w�}�Wϐ�4����t#�	N����u�u�u�<�g�
�3���D����l�N��Uʱ�;�
���w�c�D��Y���F��X��"����h�u�g�]�}�W���Ӌ��NǻN��U���9�u�k�4��1�[���Y�����R��Kʴ�
�&�y�u�w�}�WϺ������h��B���%�y�u�u�w�}����Y����A��B1�@���y�u�u�u�w�2����Y����A��B1�@���6�1�y�u�w�}�WϽ�Y����A��B1�@���y�u�u�u�w�9����GӁ��l �� \�����_�u�u�3�g�;��������]�� ��F؊�
� �9�1�'��@������]���1��a�3�e�3�3�;����K������\��*���9�1�%�u�w�:����Ӌ��NǻN��U����h�u�y�w�}�W���7����g'��S�F�ߊu�u�u�u�>�m� ���1��� T�N��U���1�;�
���}�I��U���F�
�������h�u�e�W�W�������R�=N��U���u�9�u�k�6����Y���F��R��U��4�
�&�y�w�}�W�������X��E�� ��l�%�y�u�w�}�WϺ������h��B���%�y�u�u�w�}���������h��B���:�6�1�y�w�}�W��������h��B���6�y�u�u�w�}����Y����A��B1�L���|�_�u�u�1�m����&�Ԣ�lU��D1�*ي� �9�1�%��e�MϽ�����]��\��C���3�e�3� ��o�������lU��B�����u�u�2�;�%�>����Q���F�'��H���y�u�u�u�w��:���8���F��=N��U���u�<�e����J���K���F�N��ۊ���u�k�d�q�W���Y����\��`'��=��u�g�_�u�w�2�ϳ�	��ƹF�N�����k�4�
�9�{�}�W���YӔ��V�	N��*���y�u�u�u�w�9����GӁ��l �� ]�����u�u�u�u�3�3�W�������F9��1��Y���u�u�u�6�w�c�������� 9��d��U���u�1� �u�i�:����&����CT�=d��Uʳ�e�3� �
�e�.�Dݰ�&�ԓ�l ��[1�����l�o�6�8�8�8�ϳ�K���� ��1�� ���g�&�f�;��o�D�������Cl�N�����6�8�%�}�w�}�W���0���W�N��U��������`�W��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��y�u�u�u�w�9����0����X�GךU���:�!�8�%��}�W���YӅ��[�V�����u�u�u�u�%�.���Y����@�N��U���1�;�u�k�0�-����JĹ��l�N��Uʱ�;�u�k�2�'�;�(��&����F�N�����k�2�%�3��n�(���s���F�S��U��2�%�3�
�d��E��s���U9��Q��*���&�f�;�
�e�l��������V������;�u�e��a�i�������� T��h]����
�
�4�
�$�W�W�������PF��GN��U���u�u��u�i�l�}���Y���}3��d:��0��u�y�u�u�w�}����&����{F�]����u�u�u�<�f�
�3���D����l�N��Uʱ� �
���w�c�D���Y����\��Z��]���u�u�u�1�9�}�IϹ�	����R��G^�U���u�u�1�;�w�c�������� 9��d��U���u�1� �u�i�:����&����CT�=d��Uʳ�e�3� �
�e�.�Dݰ�&�ԓ�l��h
��*��u�u�:�%�9�3�W��=����u ��h����;�
�g�&�d��(���&����F�P�����8�%�}�u�w�}�Wϗ�Y���l�N��Uʛ�����j�}�[���Y�����1��1���h�u�g�_�w�}�W����ד�z"��S�F���u�u�u�u�3�(�(���-���U��=N��U���!�8�%�}�w�}�W�������X��E�� ��m�%�y�u�w�}�WϺ������h��B���%�y�u�u�w�}����Y����A��B1�M���|�_�u�u�1�m����&�Ԣ�lU��D1�*ۊ�4�
�&�
�a�}�W���	����GF��*�Fޓ�
�
�8�9�d�3�(���
����9��O1�����u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���g�_�u�u�8�)����Q���F�
��E��u�'�
� �`�n���Y���F��^ �H���'�
� �b�d�-�[���Y�����CN��U���
� �b�f�'�t�}���YӀ��l ��[1����g�&�f�
��<�(���&����	F��Z�����8�g�e�f���(�������@9��Y��G���8�-�1�%�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�o�}���Y������FךU���u�u�<�e�j�}��������l��=N��U���u�<�d�h�w�/�(���N�ѓ�JǻN��U���:�!�h�u�%����N����lǻN��*ڊ�8�9�f�;��o���&¹��K9��G1��A��6�8�:�0�#�0�E��JǠ��9��B��G���f�;�
�g�f�0����	�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�f�W�W���Y�ƨ�]V��~*��U��f�y�u�u�w�}����&����{F�]����u�u�u�:�#�
�3���D����l�N�����4�u�_�u�w�}�W���I���U5��z;�����
� �!�%�.�l�(ށ�����l��=N��U���u�<�d�h�w�����-����l+��C����
�
� �b�f�-�[���Y�����CN��U���-� ���#���������lW��B1�D���|�_�u�u�1�m����&�Ԣ�lU��D1�*ۊ�4�
�&�
�a�}�W���	����GF��*�Fޓ�
�
�8�9�d�3�(���
����9��O1�����u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���g�_�u�u�8�)����Q���F�
��E��u��-� ����������J9��h_�� ��c�%�y�u�w�}�WϺ���� ��O#��!���!��9�<�;��C�������9��d��U���u�1� �u�i�;�(���5����G9��[�����a�d�3�
�a��E��s��ƓF�C����� �'�;�u�#�)�Wǿ�&����@�X�����!�!�u�4�?�3�Y��s���R��d1�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�4������E�ƭ�l5��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�u�w�}�W���Y���F�N�����
�&�u�h�6��$������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u�%��(߁�&�ד�F9��1��*���'�
�%�&�6�)��������]F��X�����x�u�u�2�'�;�G���H¹��lQ��h�����!�4�
�!�%�����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��G1��E���d�
� �b�a�<�(�������l��E�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����c�|�u�=�9�W�W���Y���F�N��Uʲ�%�3�e�3�f����O����@��C1��*���'�
�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}����Y�έ�l��D�����
�u�u�'���(���H����W��V�����|�u�=�;�]�}�W���Y���F�N�����3�e�3�d��(�@�������R��V�����
�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϹ�	����l ��1��*��
�%�&�4�#�<�(�������TF��D��U���6�&�{�x�]�}�W���&����U9��h��C���4�
�!�'��-��������l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�
�
�e�;�(��&����G��h�����!�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�f�3�8�f�t�^Ϫ���ƹF�N��U���u�u�u�u�%��(߁�&�ԓ�F9��1��*���'�
�%�&�6�)����E�ƭ�l��D�����
�n�u�u�w�}�W���Y����_��F�����;�!�9�2�4�l�JϹ�	����l ��1��*��
�%�'�4�.�t����Y���F�N��U���u�u�u�'���(���K����_��V�����
�%�&�4�#�/���Y����\��h�����n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��G1��E���f�3�
�a��-��������@��C1��ʴ�&�2�u�'�4�.�Y��s���T��Q1�����3�
�a�
�'�.��������R��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�2�%�1�m��������9��h�����%�&�4�!�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�c�;���PӇ����F��*���&�
�:�<��}�W���&����U9��h��C���4�
�:�0�~�t����Y���F�N��U���u�u�u�'���(���&����R��G1�����4�
�!�'��8�W������]��[����_�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����&ù�� 9��hX�*���'�4�,�|�#�8�W���Y���F�N��U���u�'�
�
���(���O�ғ�C9��V�����!�'�
�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��9��C�����0�e�4�
�;���������]F��X�����x�u�u�%�f���������V9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}���&����\��D1��E���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�w�5��ԜY���F�N��U���u�u�u�%�f���������V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�e��!�8�3����I����E
��G��U��%�d�
�0�'�4����&ù��l��d��U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�F߁�����]��R1�����u�&�<�;�'�2����Y��ƹF��h_��&���:�;�&�0�g�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��^�����<�!�
�
��/���Y����\��h��G��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	����`��X�����e�4�
�9�~�t����Y���F�N��U���u�u�u�
�g���������lV��E��I���
�e��!�8�3����I���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u��l�>�������9��h��*���2�4�&�2�w�/����W���F�G1�*��� �&�0�e�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*����%�!�
����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�}�'�>��������lW������6�0�
��$�o�(���&�����YNךU���u�u�u�u�w�}�W���Y�Ƽ�W��Y�����e�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�c�t����Y���F�N��U���u�u�u�u�w��F���	����V9��V�����'�2�i�u��l�>�������9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�H¹��C��h��*���2�4�&�2�w�/����W���F�G1�*��� �&�0�e�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��h'�� ���0�e�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(���0����@9��1��*���|�|�!�0�w�}�W���Y���F�N��U���d��%�!���(������C9��h'�� ���0�e�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���D���%�!�
�
��-����	����R��P �����&�{�x�_�w�}�(���0����@9��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�H¹��C��h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��GҊ�&�
�b�|�#�8�W���Y���F�N��U���u�u�u�
�f�����&����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��hZ�\ʡ�0�u�u�u�w�}�W���Y���F�N��*����%�!�
����������TF���D���%�!�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�d�
�;�"�.����	����R��P �����&�{�x�_�w�}�(���0����@9��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u��l�>�������9��R	��Hʴ�
�:�&�
�!�o�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���d��%�!���(������F��R ��U���u�u�u�u�w�}�W���	����z��C��*ۊ�'�2�i�u��l�>�������]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p���&����G��h\�����1�%�0�u�$�4�Ϯ�����F�=N��U���d��%�!���(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�d�
�;�"�.��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���A����lT��N�����u�u�u�u�w�}�W���Y���F��h_��<���!�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�C��Y����l�N��U���u�u�u�u�w�}�WϮ�H¹��C��h��*���#�1�%�0�w�`���&����G��h\�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�W��Y�����g�%�0�u�$�4�Ϯ�����F�=N��U���d��%�!���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���D���%�!�
�
��/���Y����\��h��G��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	����z��C��*؊�%�#�1�|�w�5��ԜY���F�N��U���u�%�d�
�9�(����K����TF���D���%�!�
�
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�d�
�;� �$�8�D���&����C�������%�:�0�&�w�p�W���	����z��C��*ي�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�W��Y�����f�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�m�3�8�e�t�W������F�N��U���u�u�u�u�w�-�Fށ�����l��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����a�u�=�;�]�}�W���Y���F�N��U���%�d�
�;�"�.��������W9��R	��Hʥ�d�
�;� �$�8�D���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
�f�����&����C�������%�:�0�&�w�p�W���	����z��C��*ي�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}���&����G��h]�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�d�
�9�(����J����E
��G�����_�u�u�u�w�}�W���Y���C9��h'�� ���0�f�%�0�w�`���&����G��h]�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����l/��B�����4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�d�
�9�(����M����E
��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
�f�����&����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���F�N����
�;� �&�2�i��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�W��Y�����a�4�
�9��/���Y����l/��B�����4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h_��<���!�
�
�
�%�:�����Ƽ�\��D@��X���u�%�d�
�9�(����M����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�d�
�;� �$�8�C��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��h'�� ���0�a�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u��l�>�������9��R	��Hʥ�d�
�;� �$�8�C�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�d��-����&ƹ��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��h'�� ���0�`�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h_��<���!�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�g��.�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&�ד�]��D1��@���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�}�W���YӃ��Z �V�����1�
�l�|�#�8�W���Y���F�N��U���u�u�u�
�f�����&����R��[
�����i�u�
�d��-����&ƹ��l��d��U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�Fށ�����l��h��ʴ�&�2�u�'�4�.�Y��s���C9��h'�� ���0�`�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����l/��B�����%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u��l�>�������9��h��\���!�0�u�u�w�}�W���Y���F���D���%�!�
�
��/���Y����l/��B�����_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����1�����
�
�
�%�!�9����Y����T��E�����x�_�u�u��l�>�������9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�Fށ�����l��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y�����T�����2�6�d�h�6�����
����g9��V�����b�|�!�0�w�}�W���Y���F�N��U���u�
�d��'�)�(���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lS��N�����u�u�u�u�w�}�W���Y���F��h_��<���!�
�
�
�'�+���������1�����
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C���
�;� �&�2�k����Y����T��E�����x�_�u�u��l�>�������9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�d��-����&Ź��V�
N��*���&�
�#�g�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���D���%�!�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}���&����G��hX�����i�u�
�d��-����&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�i�:�������G��h��*���#�1�%�0�w�.����	����@�CךU���
�
�4� �;�2����&����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�i�:�������G��h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��GҊ�&�
�b�|�#�8�W���Y���F�N��U���u�u�u�
��<��������_9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����e�|�!�0�w�}�W���Y���F�N��U���u�
�
�4�"�1��������9��h��*���2�i�u�
��<��������_9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l+��B�����:�
�
�
�%�:�����Ƽ�\��D@��X���u�%�a��9�<�4�������lV��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�a��3��������l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w��(�������]��[1��E���
�9�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\���!�0�u�u�w�}�W���Y���F���*��� �9�:�!�8��(߁����F��1������;�'�9�2�m�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�4�"�1��������9��h��*���2�4�&�2�w�/����W���F�G1��8���4��;�'�;�8�F���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�4�"�1��������9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���u�=�;�_�w�}�W���Y���F�N��Uʥ�a��;�4��3�����ד�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��_�U���;�_�u�u�w�}�W���Y���F�N��A���;�4��;�%�1��������W9��R	��Hʥ�a��;�4��3�����ד�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ہ�����p	��E�����%�0�u�&�>�3�������KǻN��*ފ�4� �9�:�#�2�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�4� �9�8�)����&¹��V�
N��*���&�
�#�g�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*��� �9�:�!�8��(ށ�	����O�C��U���u�u�u�u�w�}�W���YӖ��l+��B�����:�
�
�
�%�:�K���&ǹ��]��t�����0�d�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*��� �9�:�!�8��(݁�	����l��PN�����u�'�6�&�y�p�}���Y����~��V�����9�0�g�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*��� �9�:�!�8��(݁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����Q����ߊu�u�u�u�w�}�W���Y���F��1������;�'�9�2�o��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��Y��6���'�9�0�g�6��������F��1������;�'�9�2�o������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6�(��������V9��G��U���<�;�%�:�2�.�W��Y����lR��V �����!�:�
�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h#�� ���:�!�:�
������E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��Y��6���'�9�0�g�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(ہ�����p	��E�����%�0�u�h�'�i�:�������G��h��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Y��6���'�9�0�f�6���������@��YN�����&�u�x�u�w�-�C�������\��X��*ي�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��Y��6���'�9�0�f�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!�o�;���P�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ғ�R��[-�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�l�F������F�N��U���u�u�u�u�w�}����4����_%��C��*���
�%�#�1�'�8�W��	�ғ�R��[-�����
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����;�4��9�/����J����TF��D��U���6�&�{�x�]�}�W���&����R
��Y�����f�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ǹ��]��t�����0�f�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ہ�����p	��E�����4�
�9�|�~�)����Y���F�N��U���u�u�
�
�6�(��������V9��G��U��%�a��;�6���������l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ہ�����p	��E�����4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�a��9�<�4�������lR��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ہ�����p	��E�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���m�3�8�g�~�}����s���F�N��U���u�u�u�u�'�i�:�������G��h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�d�e�u�?�3�}���Y���F�N��U���u�u�%�a��3��������l��h�����%�0�u�h�'�i�:�������G��h��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��z�����;�'�9�0�c�-����
������T��[���_�u�u�
��<��������_9��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u����������A	��R1�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�a��3��������l��h�����|�u�=�;�]�}�W���Y���F�N������;�4��9�/����M����TF���*��� �9�:�!�8��(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�a��3��������l��h�����%�0�u�&�>�3�������KǻN��*ފ�4� �9�:�#�2�(���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�a��3��������l��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y�����T�����2�6�d�h�6�����
����g9��V�����b�|�!�0�w�}�W���Y���F�N��U���u�
�
�4�"�1��������9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��A���!�0�u�u�w�}�W���Y���F�N��U���
�4� �9�8�)����&ƹ��l��h����u�
�
�4�"�1��������9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�M����F��X �����
�
�'�2�6�.��������@H�d��Uʥ�a��;�4��3�����ӓ�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�a��;�6���������l��PN�U���6�;�!�9�d��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������;�4��9�/����L����E
��G�����_�u�u�u�w�}�W���Y���C9��z�����;�'�9�0�b�-����DӖ��l+��B�����:�
�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����;�4��9�/����O����E
��G��U���<�;�%�:�2�.�W��Y����lR��V �����!�:�
�
��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������;�4��9�/����O����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ޓ�@�� G�����u�u�u�u�w�}�W���Y���F���*��� �9�:�!�8��(ف�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������^�C��U���u�u�u�u�w�}�W���Y�����h#�� ���:�!�:�
����������TF���*��� �9�:�!�8��(ف�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�c�����:����\
��hX�����4�&�2�u�%�>���T���F��1������;�'�9�2�k����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��8���4��;�'�;�8�A��������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h#�� ���:�!�:�
���������G��d��U���u�u�u�u�w�}�WϮ�M����F��X �����
�
�'�2�k�}�(ہ�����p	��E����_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h#�� ���:�!�:�
����������TF��D��U���6�&�{�x�]�}�W���&����R
��Y�����b�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h#�� ���:�!�:�
����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�}�'�>��������lW������6�0�
��$�o�(���&�����YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��Y��6���'�9�0�b�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ǹ��]��t�����0�b�4�
�;�����E�Ƽ�9��Y��6���'�9�0�b�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�4� �;�2����&����C�������%�:�0�&�w�p�W���	�ғ�R��[-�����
�
�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l+��B�����:�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�M����F��X �����
�
�%�#�3�t�W������F�N��U���u�u�u�%�c�����:����\
��hY�����i�u�
�
�6�(��������V9��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L����T��h^�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�4�2�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�`��;�0�2�m��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�O�������F��R ��U���u�u�u�u�w�}�W���Y����lS��V ��*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�d�a�}����s���F�N��U���u�u�u�u�'�h�%�������l��A�����u�h�%�`��3����I����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(�������9��R	�����;�%�:�0�$�}�Z���YӖ��l4��P��*ڊ�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����+����l��h����u�%�6�;�#�1�D݁�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�`��;�2�8�G���&����O��_�����u�u�u�u�w�}�W���Y����a��R1��E���0�u�h�%�b���������F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(�������9��h��*���2�4�&�2�w�/����W���F�G1��'���0�0�d�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���2�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�g��.�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ƹ��]��R1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�m�|�!�2�}�W���Y���F�N��U���u�u�
�
�6�:�(���&����_��E��I���
�
�4�2���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`��3����H����TF��D��U���6�&�{�x�]�}�W���&����V9��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u������&����C��R�����:�&�
�#�e�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ߊ�4�2�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����+����l��h����u�
�
�4�0��(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`��3����K����E
��G��U���<�;�%�:�2�.�W��Y����lS��V ��*���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��e�����g�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�m�3�8�e�t�W������F�N��U���u�u�u�u�w�-�B�������lT��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��Uʥ�`��;�0�2�o��������V�
N��@���;�0�0�g�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�4�2���(���Ӈ��Z��G�����u�x�u�u�'�h�%�������l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�`��9�8����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����0�g�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u������&����C��R������;�0�0�e�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�4�2���(�������A��V�����'�6�&�{�z�W�W���&ƹ��]��R1�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ӓ�R��h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��GҊ�&�
�b�|�#�8�W���Y���F�N��U���u�u�u�
��<����&����l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��]�����u�u�u�u�w�}�W���Y���F���*���2�
�
�
�'�+���������h<�����
�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��@���;�0�0�f�'�8�W�������A	��D�X�ߊu�u�
�
�6�:�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�4�2�
������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l4��P��*ي�%�#�1�|�w�5��ԜY���F�N��U���u�%�`��9�8����	����[��h[�����
�
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��@���;�0�0�a�6���������@��YN�����&�u�x�u�w�-�B�������lR��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ځ�����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�`��;�2�8�C���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������O��_�����u�u�u�u�w�}�W���Y���C9��e�����a�4�
�9��/���Y����a��R1��A���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h<�����
�
�'�2�6�.��������@H�d��Uʥ�`��;�0�2�i����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��'���0�0�a�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����V9��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�4�2�
������E�Ƽ�9��Y	����_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h<�����
�
�%�#�3�-����
������T��[���_�u�u�
��<����&ƹ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b������ӓ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h\�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ߊ�4�2�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���H�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ӓ�R��h��*���#�1�%�0�w�`����+����l��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����a��R1��@���0�u�&�<�9�-����
���9F���*���2�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lS��V ��*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�h�%�������l��A��\���=�;�_�u�w�}�W���Y���F�G1��'���0�0�`�%�2�}�JϮ�L����T��h[�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����a��R1��C���
�9�
�'�0�<����Y����V��C�U���%�`��;�2�8�A���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�4�0��(ف�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����Q����ߊu�u�u�u�w�}�W���Y���F��1�����0�c�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ځ�����V9��V�����'�2�i�u������&����R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����+����l��h��ʴ�&�2�u�'�4�.�Y��s���C9��e�����c�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ƹ��]��R1�����u�h�4�
�8�.�(���K����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�6�:�(���&����_�N�����u�u�u�u�w�}�W���Y����lS��V ��*���
�'�2�i�w��(�������]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����+����l��h�����%�0�u�&�>�3�������KǻN��*ߊ�4�2�
�
��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������;�0�0�`�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�4��2��������F�V�����&�$��
�#�e����K���G��d��U���u�u�u�u�w�}�W���YӖ��l4��P��*݊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�g�l�w�5��ԜY���F�N��U���u�u�u�%�b������ѓ�C9��S1�����h�%�`��9�8��������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u������&����C�������%�:�0�&�w�p�W���	�ӓ�R��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�B�������lQ��E��I���%�6�;�!�;�n�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�`��;�0�2�j���������YNךU���u�u�u�u�w�}�W���&ƹ��]��R1�����u�h�%�`��3����N���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u������&����R��[
�����4�&�2�u�%�>���T���F��1�����0�m�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h[�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��@�������9F�N��U���u�u�u�u�w�}�W���&����V9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����a�|�!�0�w�}�W���Y���F�N��U���u�
�
�4�0��(ׁ�	����l��PN�U���
�4�2�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�`��9�8����	����R��P �����&�{�x�_�w�}�(ځ�����V9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��<����&˹��V�
N��*���&�
�#�g�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���2�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�B�������l^��E��I���
�
�4�2���L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�`��9�8��������W9��R	�����;�%�:�0�$�}�Z���YӖ��l4��P��*ӊ�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��Y	�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���m�3�8�g�~�}����s���F�N��U���u�u�u�u�'�h�%�������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�B���=�;�_�u�w�}�W���Y���F�N������;�0�0�n�<�(���&����Z�G1��'���0�0�l�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�4�2�
����������]F��X�����x�u�u�%�b������ߓ�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�`��;�2�8�N��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��e�����l�4�
�9�~�t����Y���F�N��U���u�u�u�
��<����&ʹ��V�
N��@���;�0�0�l�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�4�4�0�2�.��������W9��R	�����;�%�:�0�$�}�Z���YӖ��l6��V�����0�e�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hX�����0�0�&�0�g�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�4��2��������F�V�����&�$��
�#�e����K���G��d��U���u�u�u�u�w�}�W���YӖ��l6��V�����0�e�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��k�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ف�����G��h��*���#�1�%�0�w�`����)����V��D1��E���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h>�����0�&�0�e�'�8�W�������A	��D�X�ߊu�u�
�
�6�<����
����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�c��%�0����&����C��R�����:�&�
�#�e�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*܊�4�4�0�0�$�8�G���&����O��_�����u�u�u�u�w�}�W���Y����c��Z�����
�
�'�2�k�}�(ف�����G��h��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��E�����
�
�
�%�!�9����Y����T��E�����x�_�u�u����������l��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����^��E��*ۊ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�b�~�)����Y���F�N��U���u�u�u�u����������l��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����`�u�=�;�]�}�W���Y���F�N��U���%�c��'�:�)����&¹��l��h����u�
�
�4�6�8�����ד�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ف�����G��h��*���2�4�&�2�w�/����W���F�G1��%���8�!�'�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hX�����0�0�&�0�f�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����c��Z�����
�
�%�#�3�t�W������F�N��U���u�u�u�%�a���������V9��G��U��%�c��'�:�)����&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�k�'�������@9��1��*���
�'�2�4�$�:�W�������K��N������'�8�!�%��(܁�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�c��%�0����&����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���F�N������'�8�!�%��(܁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������
R�C��U���u�u�u�u�w�}�W���Y�����h>�����0�&�0�f�6��������F��1�����!�'�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�c��'�:�)����&����V��D��ʥ�:�0�&�u�z�}�WϮ�O����R��R�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����^��E��*ي�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�a���������V9��V�����|�!�0�u�w�}�W���Y���F�N��*܊�4�4�0�0�$�8�D��������h>�����0�&�0�f�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�4�;�
����������TF��D��U���6�&�{�x�]�}�W���&����@9��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�N����]��h^�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�b�|�!�2�}�W���Y���F�N��U���u�u�
�
�6�3�(���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lU��N�����u�u�u�u�w�}�W���Y���F��hY�����
�
�
�%�!�9����Y����lQ��V��*���
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��2���&�0�e�%�2�}����Ӗ��P��N����u�
�
�4�9��(߁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�4�;�
�
��/���Y����\��h��G��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ѓ�R��h��*���#�1�|�u�?�3�}���Y���F�N��U���%�b��<�$�8�G��������h)�����
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��2���&�0�d�4��1�(���Ӈ��Z��G�����u�x�u�u�'�j�0���
����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���u�=�;�_�w�}�W���Y���F�N��Uʥ�b��<�&�2�l��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��^ �����4�
�9�
�%�:�K���&Ĺ��Z��R1�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��V��*���
�'�2�4�$�:�W�������K��N������<�&�0�f�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F�� 1�����0�d�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�����V9��V�����|�!�0�u�w�}�W���Y���F�N��*݊�4�;�
�
��/���Y����t��D1��D�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��V��*���
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
�6�3�(���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�b��4����K����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ޓ�@�� G�����u�u�u�u�w�}�W���Y���F���*���;�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�D��Y����l�N��U���u�u�u�u�w�}�WϮ�N����]��h\�����1�%�0�u�j�-�@�������lT��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��Z��R1�����u�&�<�;�'�2����Y��ƹF��hY�����
�
�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l!��Y��*؊�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�`������ԓ�C9��SG��U���;�_�u�u�w�}�W���Y���F�� 1�����0�g�%�0�w�`����>����l��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��Z��R1�����9�
�'�2�6�.��������@H�d��Uʥ�b��<�&�2�n��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�4�;���(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�Eׁ�
����O��_�����u�u�u�u�w�}�W���Y���C9��p�����f�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�d�t����Y���F�N��U���u�u�u�u�w��(������� 9��h��*���2�i�u�
��<����&����l��d��U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�@�������lU��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����@9��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�4�9��(܁�	����O�C��U���u�u�u�u�w�}�W���YӖ��l!��Y��*ي�'�2�i�u������&����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�@�������lR��G1�����0�u�&�<�9�-����
���9F���*���;�
�
�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��B���<�&�0�a�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!�o�;���P�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�f�m�u�?�3�}���Y���F�N��U���u�u�%�b��4����M����E
��G��U��%�b��<�$�8�C���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��<����&ǹ��V��D��ʥ�:�0�&�u�z�}�WϮ�N����]��hZ�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�j�0���
����l��PN�U���6�;�!�9�d��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������<�&�0�c�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����@9��1�����h�%�b��>�.���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��<����&ƹ��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��p�����`�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h)�����
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��j�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*���|�!�0�u�w�}�W���Y���F�N��U���
�
�4�;���(�������A��S��*݊�4�;�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b��<�$�8�B����ƭ�@�������{�x�_�u�w��(�������9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�6�3�(���&����Z�V�����
�#�g�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY�����
�
�
�%�!�9�^������F�N��U���u�u�u�u�'�j�0���
����l��PN�U���
�4�;�
��f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b��<�$�8�A���&����C�������%�:�0�&�w�p�W���	�ѓ�R��h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����t��D1��C���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�w�5��ԜY���F�N��U���u�u�u�%�`������Г�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��X�U���;�_�u�u�w�}�W���Y���F�N��B���<�&�0�c�6��������F�� 1�����0�c�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��/�Ͽ�
����C��R��U���u�u�%�b��4����O����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��<�&�2�k����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��^ �����4�
�9�|�~�)����Y���F�N��U���u�u�
�
�6�3�(���&����Z�G1��2���&�0�c�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*݊�4�;�
�
��-����	����R��P �����&�{�x�_�w�}�(؁�����V9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����>����l��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y�����T�����2�6�d�h�6�����
����g9��V�����b�|�!�0�w�}�W���Y���F�N��U���u�
�
�4�9��(؁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������S�C��U���u�u�u�u�w�}�W���Y�����h)�����
�
�%�#�3�-����DӖ��l!��Y��*݊�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�����0�b�%�0�w�.����	����@�CךU���
�
�4�;���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���;�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N����]��hY�����1�|�u�=�9�W�W���Y���F�N��Uʥ�b��<�&�2�j����Y����lQ��V��*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�����0�m�4�
�;���������]F��X�����x�u�u�%�`������ޓ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u������&����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���F�N������<�&�0�o�<�(���&����Z�V�����
�:�<�
�l�}�W���Y���F�N��U���<�u�4�
�>�����A����[��=N��U���u�u�u�u�w�}�W���Y����t��D1��M���
�9�
�'�0�a�W���&����@9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l!��Y��*Ҋ�'�2�4�&�0�}����
���l�N��B���<�&�0�m�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��p�����m�%�0�u�j�<�(���
���� T��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������9��h��\���!�0�u�u�w�}�W���Y���F���*���;�
�
�
�%�:�K���&Ĺ��Z��R1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ӊ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�4�9��(ց�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�b��>�.��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���A����lT��N�����u�u�u�u�w�}�W���Y���F��hY�����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�n�D������F�N��U���u�u�u�u�w�}����>����l��h�����%�0�u�h�'�j�0���
����l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����@9��1�����&�<�;�%�8�8����T�����h)�����
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ѓ�R��h��*���2�i�u�%�4�3����J����9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�b��4����@����E
��G�����_�u�u�u�w�}�W���Y���C9��p�����l�%�0�u�j�-�@�������l_��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R
��R1�����9�
�'�2�6�.��������@H�d��Uʥ�l��2�4�$�8�G���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�<�9�1�(���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���K˹��^9��G�����_�u�u�u�w�}�W���Y���F�G1��&���4�&�0�e�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ʹ��T��D1��E���
�9�
�'�0�a�W���&����R
��R1�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����l_��^	�����
�
�'�2�6�.��������@H�d��Uʥ�l��2�4�$�8�G�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��L���2�4�&�0�g�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l5��Y��*���
�%�#�1�~�}����s���F�N��U���u�u�%�l��:�����֓�A��S��*ӊ�<�;�9�
��f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�l��2�6�.��������W9��R	�����;�%�:�0�$�}�Z���YӖ��l5��Y��*���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��d�����0�d�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�m�3�:�o�^������F�N��U���u�u�u�u�w�}����*����_��h_�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����a�d�u�=�9�W�W���Y���F�N��U���u�%�l��0�<����H����E
��G��U��%�l��2�6�.��������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������9��R	�����;�%�:�0�$�}�Z���YӖ��l5��Y��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�@����]��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��4����&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��hW�����9�
�
�
�%�:�K���&ʹ��T��D1��D�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����l_��^	�����
�
�%�#�3�-����
������T��[���_�u�u�
��4����&����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�d�$�������lT��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�<�;�;��(݁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������V�C��U���u�u�u�u�w�}�W���Y�����h=�����
�
�
�%�!�9����Y����l_��^	�����
�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��L���2�4�&�0�e�-����
������T��[���_�u�u�
��4����&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�<�9�1�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��&���4�&�0�g�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(ց�����@9��1�����h�%�l��0�<����K���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��Z�����f�u�;�u�8�u��������_	��T1�Hʲ�%�3�e�3�f����@����W	��G��U���;�u�u�u�w�}�W���YӅ��u#��u/����� �
�l�e�2�m�K�������9��\�� ��l�4�
�0�"�3�G�ԜY���F�N��Uʶ�
�:�0�!�%�����)����c*��D��D���2�d�m�u�j�:����I����9��hX�*���'�!�'�
�l�}�W���Y���F������
�0�8��%�8����)����A��h��*��d�i�u�'���(���K����_��V�����;�g�_�u�w�}�W���Y���U5��X
�����
�=�0��6�8�;�������T9��X��Hʲ�%�3�e�3�f����@����A��E ��N���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B���F������%�:�0�&�w�p�W���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&�����Yd��U���u�u�u�u�w�>�(���=����\��B��L���e�'�2�d�f�}�JϽ�&����q'��X�� ���l�e�0�e�]�}�W���Y���F�Q=��&����!�d�
��8�(��A���T��Q��Fي�g�_�u�u�w�}�W���Y�ƪ�l��u����
�
�0�
�`�n�K�������lQ��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���R��Y��]���6�;�!�9�0�>�G������lV��h]�� ��a�4�
�:�2�t�^Ϫ����F�N��U���u�6�
�:�2�)��������V��Y�����d�'�2�d�g�}�JϹ�	����l ��h��C���4�
�0� �9�l�}���Y���F�N�����:�0�!�'��<��������A	��D1�����d�d�u�h�0�-�����Փ�F9��1��*��� �;�g�_�w�}�W���Y���F��h �����'�
�4�6�3�9�������� 9��P1�D���h�2�%�3�g�;�D���&����R��R����_�u�u�u�w�}�W���Y����\��C��*���6�1�1�:�#�2�(���&����^��R�����3�e�3�f�1��Cہ�	����F��UךU���u�u�u�u�w�}��������A��V�����:�!�:�
������A���F��G1��E���f�3�
�a��-��������9F�N��U���u�u�u�9�9�9�(�������P��S-�����
�
�
�0��e�E��Y����U9��Q1�����a�
�%�'�#�/�(��Y���F�N��U���9�;�1�
�2�0�4�������\��X��*݊�0�
�m�b�k�}����&ù�� 9��hX�*���'�!�'�
�l�}�W���Y���F������
�0�8��$�<��������l��h��*��g�i�u�'���(���&����R��G1�����
�n�u�u�w�}�W���Y����_9��S������&�4�0��3����
�ߓ�V��Z�I���'�
�
�
�����M����A��E ��N���u�u�u�u�w�}�WϽ�&����l��Z1�����0��;�'�;�.����H����[��E��*ڊ�
�
� �c�c�<�(�������l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�e�3�:�l�^�������F�N��U���u�u�3�
���#���&�Г�l��h_�E��u��������&����lW��1��N���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B���F������%�:�0�&�w�p�W���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�@�������O��_��U���u�u�u�u�w�}����<����|��^��*���
�m�a�i�w��$���:����l^��1��*��l�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U�� G�����:�}�4�
�8�.�(�������F��G1��E���d�
� �b�a�<�(��������Yd��U���u�u�u�u�w�;�(�������^9��Y��&���<�g�
�0��j�O��Y����U9��Q1�*���b�c�4�
�2�(���s���F�N��U���3�
�:�0�#�/�(���������_�����b�a�i�u�%��(߁�&�ד�F9��1��*��� �;�d�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-���� 9��Z1�\���!�0�_�u�w�}�W���Y���U5��v*��:���g�
�
�0��j�E��Y����U��[��G�ߊu�u�u�u�w�}�W���*����q��C1�����6�
�m�d�%�:�F��Y����A��B1�L���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����VO��Y
�����%�&�2�7�3�j�@���Y����9F�N��U���u�u�u��/��#ݰ�����lW��R	��B��i�u��-��	����&�֓�l ��^�*��_�u�u�u�w�}�W���Y����~3�� ����
�
�0�
�`�k�K���*����2��x��Gڊ�
� �d�l��n�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�6�.��������@H�d��Uʥ�:�0�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��|�!�0�_�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����g�|�|�!�2�W�W���Y���F�N��*����g��!�`�l����H����[��d1�� ���;� �
�
��(�F��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�t�W������F�N��U���u��-� ����������J9��h_�����b�b�i�u�%����A����9F�N��U���u�u�u��/��#�������G��N1�*ۊ�0�
�b�b�k�}��������l��=N��U���u�u�u�u�w�����-����l+��C�����d�'�2�d�a�}�JϹ�	����S��G\�U���u�u�u�u�w�}����4����|��z�����
�
�
�0��j�E��Y����U��]��G�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�N������F��R ךU���u�u�u�u�w�}�$���,����F��B�����d�
�
�0��j�A��Y����~3��N!��*���!�%�,�d�����O����9F�N��U���u�u�u��/��#�������G��N1�*ۊ�0�
�b�e�k�}�$���,����F��B�����d�
�
� �`�l���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Gފ�&�
�f�|�w�5����Y���F�N��U���-� �,� ������A���F��G1��*��
�g�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�b�3�8�a�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��_��\���=�;�u�u�w�}�W���Y����V�� ]��Hʲ�%�3�
�g��o�}���Y���F�N�����b�d�i�u�%����@����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����T��E�����x�_�u�u�%�>��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�r�p�}����Y���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�������R��X ��*���<�
�u�u�%��(߁�&�ד�F9��1��*���0�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&���\������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�u�;�w�2�_ǿ�&����G9��P��E��2�%�3�e�1�l�(���O�ߓ�C9��Y��U���u�:�}�4��2����¹��F��1�����&�0�g�'�6���������9��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��m�^ϱ�Y�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���u�=�;�u�w�}�W���Y�����hY�U��2�%�3�
�c��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��M���8�b�u�;�w�2�_ǿ�&����G9��P��E��2�%�3�e�1�l�(���N�Г�C9��Y��\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�l�3�:�e�^ϱ�Y�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\ʴ�1�;�!�}�'�>��������lV�	��*���
�
�g�3��d�(�������F��SN�����%�6�;�!�;�l�G��	�ߓ�Z��[��*؊�0�1�'�4��(�E���	���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��D���8�g�|�|�w�5����Y���F�N��U���
�l�u�h�0�-����M˹��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�l�3�:�e�^ϱ�Y�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���u�=�;�u�w�}�W���Y�����hV�U��2�%�3�
�b��E�ԜY���F�N��Uʧ�2�m�l�i�w�/�(���N�ѓ�]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�4�
�8�.�(�������F��h��U���u�:�}�4��2����¹��F��1�����&�0�g�'�6���������9��G�����4�
�:�&��2����Y�ƭ�l��h�����
�!�b�3�:�l�^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����R��D��F���|�!�0�_�w�}�W���Y���F��P1�A��u�'�
� �`�d���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}��������G��F��*���3�8�u�3�#�8����Ӌ��[��N����u�%��
�$���������PF��G�����}�%��
�$�q�����ƫ�C9��1��Dۊ� �b�c�4��2��������9��\�� ��l�4�
�:�2�}��������lQ��N�����e�3�f�3��i�(�������9F����ߊu�u�u�u�6�8����*������N��U���u�u�"�0�w�-�$���¹��^9��
P��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�����έ�l��h��*��|�|�!�0�]�}�W���Y���F�N������3�8�i�w�-�$�������^9��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��D��N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�-�9���
�����d:��ي�&�
�n�u�w�}�W���Yӑ��]F��h=�����3�8�g�h�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�"�0�u�'��(���&���� F�d��U���u�u�u�u�w�<�(������F��h=�����3�8�a�_�w�}�W���Y�ƻ�V��G1��*���
�&�
�u�i�W�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�=�;�6��#���O����lS�	NךU���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y����[��V��!���b�3�8�c�j�}�W���Y���F�N�����
�&�u�h�6��#���A����lQ��N��U���u�u�"�0�w�-�$���˹��^9��
P��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������C9��Y�����6�e�h�2�'�;�G���H¹��lQ��h�����|�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
�ߓ�@��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��B�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���&����F�d��U���u�u�u�u�w�<�(������F��h=����
�&�
�n�w�}�W���Y����[��V��!���d�
�&�
�w�c�}���Y���F�N������3�8�i�w�-�$����ד�@��UךU���u�u�u�u�?�3����-����9��Z1�U��_�u�u�u�w�}�W���Y����`9��ZN�U����
�!�g�1�0�F��Y���F�N�����4�
��&�f�����H���9F�N��U���u�u�u�%������DӇ��`2��C_�����d�n�u�u�w�}�W�������R��c1��Dي�&�
�g�h�w�}�W���Y���F���;���&�u�h�4��	���&����U��N��U���u�u�"�0�w�-�$����ғ�@��N��U���u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y������T�����2�6�e�h�0�-��������U��W�����;�|�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�
���F�N��U���u�u�u�4������E�ƭ�l5��D�*���
�f�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����S��D��A��u�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	�������!�9�2�6�g�`�����֓�lU��B1�A���
�:�0�|�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*���_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�d�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��1����u�k�_�u�w�}�W���Y���R��d1����u�%��
�#�j����H��ƹF�N��U���=�;�4�
��.�F؁�
����[�=N��U���u�u�u�u�w�-�9���
�����d:�����3�8�d�n�w�}�W���Y����[��V��!���d�
�&�
�`�`�W���Y���F�N��U����
�&�u�j�<�(���
����U��V�U���u�u�u�u� �8�W���*����_��D��M��u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�g��.�(��s���F�N�����u�%��
�#�m����H���l�N��U���u�u�u�4������E�ƭ�l5��D�*���
�e�_�u�w�}�W���Y������d:�����3�8�g�u�i�W�W���Y���F�N��*���3�8�i�u�'��(���K����lT��=N��U���u�u�u�=�9�<�(���
����U��_��K�ߊu�u�u�u�w�}�W���	����U��S�����
�!�f�3�:�o�L���Y���F���ʴ�
��&�g��.�(��D��ƹF�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�f�h�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Eځ�
����l�N��U���u�"�0�u�'��(���L����lT��
P��U���u�u�u�u�w�}����*����Z�V��!���g�
�&�
�b�W�W���Y���F��R �����
�!�c�3�:�o�W���s���F�N��U���4�
��3�:�a�W���*����Q��D��C�ߊu�u�u�u�w�}��������l�� 1����u�k�_�u�w�}�W���Y���R��d1����u�%��
�#�e����K��ƹF�N��U���=�;�4�
��.�Eׁ�
����[�=N��U���u�u�u�u�w�-�9���
�����d:��ۊ�&�
�n�u�w�}�W���Yӑ��]F��_��U��u�u�u�u�w�}�W���YӇ��}5��D��H���������/���!����k>��o6�����u�u�u�;�w�<��ԜY�Ʃ�WF��X���ߠu�u�x�u�'�9����
������T��[���_�u�u�%�3�3�(�������A	��N�����&�4�
�0�w�-��������`2��C\�����g�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��GҊ�&�
�b�|�w�5��ԜY���F�N��*���0�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������]�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����^
��U���<�;�%�:�2�.�W��Y����C9��[�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&��ƹF��R	�����u�u�u�3��3����	����@��X	��*���u�%�&�4�#�t����Q����\��h�����u�u�%�&�0�>����-����l ��h^��\ʡ�0�u�u�u�w�}�W�������_�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�>�1�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������@��YN�����&�u�x�u�w�<�(�������@��h����%�:�0�&�6�����	����l��F1��*���m�3�8�g�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��j�^������F�N��U���4�
�0�1�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�7�1�f�i�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(�������]��[1��E���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�C��Y�έ�l��D�����
�u�u�
��<��������_9��1��*���|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�G�U���0�1�%�:�2�.�}�ԜY�����D�����d�`�u�&�>�3�������KǻN�����2�7�1�d�b���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����I���F��G1�����9�d�d�h�6��$�������W	��C��B���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�e�b�<����Y����V��C�U���4�
�<�
�3��G�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������P��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�f�j�W�������A	��D�X�ߊu�u�%�&�0�?���N����@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9�� \��H���%�6�;�!�;�l�F������l ��Z�����:�a�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��G������]F��X�����x�u�u�4��4�(���&����l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�L��u�4�
�:�$��ށ�Y�ƭ�l%��Q��D���:�;�:�d�~�f�W�������A	��D����u�x�u�%�$�:����H����R��P �����&�{�x�_�w�}��������lW��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����m�u�h�}�'�>�����ד�[��G1��*���}�b�1�"�#�}�@���s���V��G�����_�_�u�u�z�<�(���&����V�������%�:�0�&�w�p�W�������T9��S1�Lي�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�e�f�k�}��������_��N������3�8�g�w�2����K���9F���U���6�&�n�_�w�}�Z���	����l��h_�U���<�;�%�:�2�.�W��Y����C9��P1����f�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��A���;�4��;�%�1��������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��D���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ǹ��]��t�����0�d�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��Y��6���'�9�0�g�6�����Y����V��=N��U���u�u�u�u�w�-��������T�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u����������A	��R1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�l�FϿ�
����C��R��U���u�u�4�
�>�����J¹��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ہ�����p	��E�����4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�F��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�4� �;�2����&����R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�d�e�4�$�:�W�������K��N�����<�
�1�
�c���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�6�(��������V9��V�����u�u�7�2�9�}�W���Y���F������7�1�d�e�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hZ�����9�:�!�:���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Lʴ�&�2�u�'�4�.�Y��s���R��^	�����a�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ފ�4� �9�:�#�2�(���&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��D��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ғ�R��[-�����
�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��V�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lR��V �����!�:�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����S��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�i�:�������G��h��*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��B������]F��X�����x�u�u�4��4�(���&����l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�G��u�4�
�:�$��ށ�Y�ƭ�l%��Q��@ʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@�ƭ�@�������{�x�_�u�w�-��������_��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��D��u�h�}�%�4�3����H�����t=�����`�1�"�!�w�h�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������R��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��X�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�c�a�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��Y�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��8���4��;�'�;�8�@���&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R
��Y�����b�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����H����@��YN�����&�u�x�u�w�<�(���&����Q��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����a��R1��E���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�A��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�4�2�
����������F�R �����0�&�_�_�w�}�ZϿ�&����Q��V����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���2�
�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�b������ד�C9��SG����u�;�u�'�4�.�L�ԶY���F��h��*���
�l�u�&�>�3�������KǻN�����2�7�1�d�c�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�`��9�8��������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��L���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ƹ��]��R1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�o�DϿ�
����C��R��U���u�u�4�
�>�����I����@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ځ�����V9��V�����u�u�7�2�9�}�W���Y���F������7�1�g�f�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h[�����
�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��\�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lS��V ��*���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�`��;�2�8�C���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��G���&�<�;�%�8�8����T�����D�����g�d�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^�����;�0�0�b�<�(���P�����^ ךU���u�u�u�u�w�}��������lT��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������9��h��\��u�u�0�1�'�2����s���F������7�1�g�e�6�.��������@H�d��Uʴ�
�<�
�1��n�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��<����&Ź��l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����e�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l4��P��*܊�%�#�1�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ϯ�L����T��hY�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�d�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��@���;�0�0�b�6�����B����������n�_�u�u�z�}��������lT�������%�:�0�&�w�p�W�������T9��S1�M���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����0�m�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����K���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�6�:�(���&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����b�4�&�2�w�/����W���F�V�����1�
�`�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�4�2���(������F�U�����u�u�u�u�w�}�WϿ�&����Q��[�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����+����l��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�a�}����Ӗ��P��N����u�%�&�2�5�9�E�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�k�'�������@9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�g�a�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���4�0�0�&�2�m�������9F���U���6�&�n�_�w�}�Z���	����l��h\�U���<�;�%�:�2�.�W��Y����C9��P1����`�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��C���'�8�!�'���(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Y�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����)����V��D1��D���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����^��E��*ي�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��N���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�c��'�8�#�/�(���&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����g�4�&�2�w�/����W���F�V�����1�
�d�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�4�;���(������F�U�����u�u�u�u�w�}�WϿ�&����Q��_�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����>����l��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�e�}����Ӗ��P��N����u�%�&�2�5�9�D�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�j�0���
����l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�g�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��p�����d�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����J����@��YN�����&�u�x�u�w�<�(���&���� U��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����t��D1��G���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�n�G��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�4�;�
����������F�R �����0�&�_�_�w�}�ZϿ�&����Q��]����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���;�
�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������
F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�`������Փ�C9��SG����u�;�u�'�4�.�L�ԶY���F��h��*���
�a�u�&�>�3�������KǻN�����2�7�1�f�o�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�b��>�.��������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��A���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��Z��R1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�n�@Ͽ�
����C��R��U���u�u�4�
�>�����LĹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(؁�����V9��V�����u�u�7�2�9�}�W���Y���F������7�1�f�b�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY�����
�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��X�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lQ��V��*���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�b��<�$�8�A���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��B���&�<�;�%�8�8����T�����D�����f�`�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^�����<�&�0�`�<�(���P�����^ ךU���u�u�u�u�w�}��������lU��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������9��h��\��u�u�0�1�'�2����s���F������7�1�f�a�6�.��������@H�d��Uʴ�
�<�
�1��e�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��<����&˹��l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����a�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l!��Y��*Ҋ�%�#�1�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ϯ�N����]��hW�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�n�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��B���<�&�0�l�6�����B����������n�_�u�u�z�}��������lR�������%�:�0�&�w�p�W�������T9��S1�G���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����&�0�e�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��4����&����R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�a�d�4�$�:�W�������K��N�����<�
�1�
�f���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�>�3����&¹��l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����d�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l5��Y��*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����K�ƭ�@�������{�x�_�u�w�-��������V��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ߓ�Z��[��*؊�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��E���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�l��2�4�$�8�E���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��G���&�<�;�%�8�8����T�����D�����a�l�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^���
�0�%�<�#��(߁�	����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�Hù��G��Y�����4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Z��H���%��
�&��}�������F��h�����#�
�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��C���
������T��[���_�u�u�%�$�:����M�ѓ�@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q���&����G��h^�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�c�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��Dۊ�;� �&�0�g�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��X�����;�%�:�0�$�}�Z���YӇ��@��U
��A���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�*��� �&�0�d�6�����Y����V��=N��U���u�u�u�u�w�-��������P�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u��l�>�������9��h��\��u�u�0�1�'�2����s���F������7�1�a�`�6�.��������@H�d��Uʴ�
�<�
�1��k�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
�f�����&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����a�`�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lW��~ �����
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lR��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��9��G��*���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�d�
�;�"�.��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�a�f�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�d�
�;� �$�8�C���&����9F����ߊu�u�u�u�w�}�W���	����l��hZ�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���H����F��R1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�i�EϿ�
����C��R��U���u�u�4�
�>�����@����@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(���0����@9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�a�e�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���D���%�!�
�
��-����P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Eۊ�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��h_��<���!�
�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�f�����
����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�d�u�$�4�Ϯ�����F�=N��U���&�2�7�1�b�o��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����L���F��G1�����9�d�d�h�6��$�������\��XN�\�ߊu�u�;�u�%�>���s���K�V�����1�
�g�u�$�4�Ϯ�����F�=N��U���&�2�7�1�b�l��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����L���F��G1�����9�d�d�h�6��$�������\��XN�\�ߊu�u�;�u�%�>���s���K�V�����1�
�f�u�$�4�Ϯ�����F�=N��U���&�2�7�1�b�m��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����L���F��G1�����9�d�d�h�6��$�������W	��C��D���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�a�w�.����	����@�CךU���%�&�2�7�3�h�D���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(��������Y��B���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�`�w�.����	����@�CךU���%�&�2�7�3�h�B���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(��������Y��M���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�c�w�.����	����@�CךU���%�&�2�7�3�h�C���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(������ F��@ ��U��|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�o�}����Ӗ��P��N����u�%�&�2�5�9�B�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������W�
N�����;�!�9�d�f�`����*����T��S�����e�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��d�W�������A	��D�X�ߊu�u�%�&�0�?���I����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lS��R��]���6�;�!�9�f�l�JϿ�&����@�N�����u�a�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��G���
������T��[���_�u�u�%�$�:����O�ѓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��Y��H���%�6�;�!�;�l�F������l ��_����!�u�c�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��hX�U��}�%�6�;�#�1�F��DӇ��p5��D��Fʱ�"�!�u�f�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����I�ƭ�@�������{�x�_�u�w�-��������Q��D�����:�u�u�'�4�.�_���
����F��1������;�'�9�2�m��������l��N��A���;�4��;�%�1��������W9��h��Yʥ�a��;�4��3�����ԓ�C9��S1��*���y�%�a��9�<�4�������lU��G1�����
�<�y�%�c�����:����\
��hZ�����1�<�
�<�{�-�C�������\��X��*ߊ�%�#�1�<��4�[Ϯ�M����F��X �����
�
�%�#�3�4�(���UӖ��l+��B�����:�
�
�
�'�+����&������h<�����
�
�%�#�3�4�(���UӖ��l4��P��*ۊ�%�#�1�<��4�[Ϯ�L����T��h\�����1�<�
�<�{�-�B�������lU��G1�����
�<�y�%�b������ғ�C9��S1��*���y�%�`��9�8��������W9��h��Yʥ�`��;�0�2�k��������l��N��@���;�0�0�b�6���������F��1�����0�m�4�
�;������Ƽ�9��Y	�����4�
�9�
�9�.����&Ź��A��C��*���
�%�#�1�>����	�Г�R��R�����d�4�
�9��3����Y����c��Z�����
�
�%�#�3�4�(���UӖ��l!��Y��*ڊ�%�#�1�<��4�[Ϯ�N����]��h_�����1�<�
�<�{�-�@�������lT��G1�����
�<�y�%�`������Փ�C9��S1��*���y�%�b��>�.��������W9��h��Yʥ�b��<�&�2�h��������l��N��B���<�&�0�c�6���������F�� 1�����0�b�4�
�;������Ƽ�9��^ �����4�
�9�
�9�.����&Ĺ��Z��R1�����9�
�;�&�0�}�(ց�����@9��1��*���
�;�&�2�w��(�������V9��V�����;�&�2�u����������9��h��*���&�2�u�
�g���������lV��G1�����
�<�y�%�f�����
����l��A�����<�y�%�d��3�����ד�C9��S1��*���y�%�d�
�9�(����K����E
��^ �����%�d�
�;�"�.��������W9��h��Yʥ�d�
�;� �$�8�C���&����Z��^	���
�;� �&�2�h��������l��N��Dۊ�;� �&�0�a�<�(���&����Z�N�����;�u�u�u�w�}�W���YӇ��@��U
��B��i�u�}�
�f�����&����R��[
�����2�h�4�
�8�.�(�������	����D���%�!�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�H¹��C��h��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�d�
�9�(����J����E
��^ �����u�%�6�;�#�1����I�ƣ�N��_�����&�0�g�4��1�(���
�����T�����2�6�e�u�%�u�(���0����@9��1��*���
�;�&�2�j�<�(���
����T��G�����
�d��%�#��(߁�	����l��D��Hʴ�
�:�&�
�8�4�(�������lW��d�����&�0�e�4��1�(���
�����T�����2�6�e�u�%�u�(ց�����@9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�<�;�;��(ށ�	����l��D��Hʴ�
�:�&�
�8�4�(�������l_��^	�����
�
�%�#�3�4�(���Y�ƭ�l��D�����
�|�:�u�'�j�0���
����l��A�����<�u�u�%�4�3��������F��F��B���<�&�0�m�6���������[��G1�����9�2�6�e�w�/�_���&����@9�� 1��*���
�;�&�2�j�<�(���
����T��G�����
�
�4�;���(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l!��Y��*ߊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�b��4����M����E
��^ �����u�%�6�;�#�1����I�ƣ�N�� 1�����0�f�4�
�;���������C9��Y�����6�e�u�'���(�������9��h��*���&�2�h�4��2��������O��EN��*݊�4�;�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�N����]��h^�����1�<�
�<�w�}��������\��h^�����%�c��'�:�)����&����l��h�����h�4�
�:�$�����&����AF��hX�����0�0�&�0�f�<�(���&����Z������!�9�2�6�g�}����&Ź��A��C��*���
�%�#�1�>�����Y����\��h�����|�:�u�%�b������ߓ�C9��S1��*���u�u�%�6�9�)�������\�G1��'���0�0�m�4��1�(���
�����T�����2�6�e�u�%�u�(ځ�����V9��V�����;�&�2�h�6�����&����P9����]���
�4�2�
����������@��
N��*���&�
�:�<��t����	�ӓ�R��h��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�`��9�8��������W9��h��U���%�6�;�!�;�:���Y���C9��e�����f�4�
�9��3����DӇ��P	��C1�����e�u�'�}������&����R��[
�����2�h�4�
�8�.�(�������	����*���2�
�
�
�'�+����&����F��h�����:�<�
�|�8�}����+����l��h�����<�
�<�u�w�-��������Z��N��U¥�a��;�4��3�����ѓ�C9��S1��*���u�u�%�6�9�)�������\�G1��8���4��;�'�;�8�A���&����Z��^	��U���6�;�!�9�0�>�G����μ�9��Y��6���'�9�0�`�6���������[��G1�����9�2�6�e�w�/�_���&����R
��Y�����a�4�
�9��3����DӇ��P	��C1�����e�u�'�}����������A	��R1�����9�
�;�&�0�`��������_	��T1�U���}�
�
�4�"�1��������9��h��*���&�2�h�4��2��������O��EN��*ފ�4� �9�:�#�2�(���&����_��Y1����4�
�:�&��2����PӉ����h#�� ���:�!�:�
����������@��
N��*���&�
�:�<��t��������R��
N��*���&�
�:�<��t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����g�i�u�4��2����¹��F��h-�����l�1�"�!�w�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����a�i�u�4��2����¹��F��h-�����d�u�:�;�8�l�^��Y����]��E����_�u�u�x�w�-��������W��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��Z�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����m�d�i�u�6�����&����F�V��&���8�d�u�:�9�2�F���B����������n�_�u�u�z�}��������l^�������%�:�0�&�w�p�W�������T9��S1�@���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�m�`�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��V�����;�%�:�0�$�}�Z���YӇ��@��U
��M���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�m�m�k�}��������_��N������3�8�g�w�2����K���9F���U���6�&�n�_�w�}�Z���	����l��F1��*���e�3�8�l�6�.��������@H�d��Uʴ�
�<�
�&�&��(���I����l_��D�����:�u�u�'�4�.�_���
����W��\��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��M��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�e�3�:�d�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�l�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�d�3�8�f�}����Ӗ��P��N����u�%�&�2�4�8�(���
����U��^�����;�%�:�u�w�/����Q����Z��S
��E��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�e�l�u�?�3�}���Y���F�V�����&�$��
�#�l����H�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$����ד�@��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�o����H�ƭ�@�������{�x�_�u�w�-��������`2��C_�����d�
�&�<�9�-����Y����V��V�����1�
�f�|�w�}�������F���]���&�2�7�1�b�m�W������F�N��Uʴ�
�<�
�&�&��(���K����lW��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���J����lW��V�����'�6�&�{�z�W�W���	����l��F1��*���f�3�8�d��.����	����	F��X��´�
�<�
�1��o�^���Yӄ��ZǻN��U���3�}�%�&�0�?���M�Ƹ�V�N��U���u�u�4�
�>�����*����U��D��G��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��Dي�&�
�g�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�>�����*����R��D��Fʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�a�1�0�F܁�
����l��TN����0�&�4�
�>�����O��ƹF��R	�����u�u�u�3��-��������R�C��U���u�u�u�u�w�<�(���&����l5��D�*���
�f�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��n�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�*���
�a�4�&�0�}����
���l�N��*���
�&�$���)�B�������R��P �����o�%�:�0�$�<�(���&����R��=N��U���<�_�u�u�w�}����	����l��hV�\ʡ�0�u�u�u�w�}�W�������T9��R��!���d�
�&�
�c�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�f�����M���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���d�
�&�
�b�<����Y����V��C�U���4�
�<�
�$�,�$����Г�@��1�����
�'�6�o�'�2��������T9��S1�L���u�u�7�2�9�}�W���Yӏ����D�����d�l�|�!�2�}�W���Y���F��G1�����0�
��&�f�����L���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���HŹ��^9��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�����OӇ��Z��G�����u�x�u�u�6�����
����g9��Y�����c�4�&�2��/���	����@��G1�����1�c�b�_�w�}����s���F�^�����<�
�1�
�g�t����Y���F�N��U���&�2�6�0��	���&����P�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����GW��Q��D���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	���&����Q��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=����
�&�
�b�6�.���������T��]���&�2�7�1�f�e�^���Yӄ��ZǻN��U���3�}�%�&�0�?���A����[��=N��U���u�u�u�%�$�:����&����GW��Q��D���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GW��Q��D���&�<�;�%�8�8����T�����D�����
��&�d��.�(�������]9��X��U���6�&�}�%�$�:����H����9F����ߊu�u�u�u�1�u��������lW��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�l�1�0�F���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ۊ�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�F����֓�@��Y1�����u�'�6�&��-��������OǻN�����_�u�u�u�w�;�_���
����W��G�����_�u�u�u�w�}�W���
����@��d:��ۊ�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C\�����d�u�&�<�9�-����
���9F������6�0�
��$�o�(���&�ߓ�@��Y1�����u�'�6�&��-��������S�N�����;�u�u�u�w�4�Wǿ�&����Q��Y�U���;�_�u�u�w�}�W���	����l��F1��*���e�3�8�d�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!�g�;���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���d�3�8�g�w�.����	����@�CךU���%�&�2�6�2��#���K¹��^9��h�����%�:�u�u�%�>����	����l��h[�\���u�7�2�;�w�}�W�������C9��P1�����d�u�=�;�]�}�W���Y���R��^	������
�!�d�1�0�E���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$����������F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�g�1�0�E���
������T��[���_�u�u�%�$�:����&����GT��Q��Gۊ�&�<�;�%�8�}�W�������R��^	�����e�f�_�u�w�8��ԜY���F��F��*���
�1�
�e�d�}����s���F�N�����<�
�&�$����������F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����T��D��D��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���������� F��D��U���6�&�{�x�]�}�W���
����@��d:�����3�8�g�
�$�4��������C��R�����<�
�1�
�f�t�W�������9F�N��U���}�%�&�2�5�9�A��Y����l�N��U���u�4�
�<��.����&����l ��h\�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(���&����l5��D�*���
�f�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��.����&����l ��h\����2�u�'�6�$�s�Z�ԜY�ƭ�l��h�����
�!�`�3�:�o�(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��[�����a�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���g�
�&�
�c�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9��X�����`�4�&�2�w�/����W���F�V�����&�$��
�#�k����Kƹ��@��h����%�:�0�&�6���������OǻN�����_�u�u�u�w�;�_���
����W��V�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�`�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�g��.�(��E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�b�6�.��������@H�d��Uʴ�
�<�
�&�&��(���A����lT��V�����'�6�o�%�8�8�ǿ�&����Q��^�\���u�7�2�;�w�}�W�������C9��P1����`�|�!�0�w�}�W���Y�����D�����
��&�g��.�(��E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	���&����Q�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�g�1�0�FϿ�
����C��R��U���u�u�4�
�>�����*����9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��D��|�u�u�7�0�3�W���Y����UF��G1�����1�d�c�|�#�8�W���Y���F������6�0�
��$�o����H���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���K����lW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�a�1�0�DϿ�
����C��R��U���u�u�4�
�>�����*����9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��@��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�d�|�!�2�}�W���Y���F��G1�����0�
��&�c�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�`�3�:�i�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�B���u�u�7�2�9�}�W���Yӏ����D�����d�b�|�!�2�}�W���Y���F��G1�����0�
��&�b�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�c�3�:�h�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�M���u�u�7�2�9�}�W���Yӏ����D�����d�m�|�!�2�}�W���Y���F��G1�����0�
��&�a�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�b�3�:�k�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�D�ߊu�u�0�<�]�}�W���Y���R��^	�����g�|�!�0�w�}�W���Y�����D�����
��&�b�1�0�A��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�@������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�m�3�8�`�<����Y����V��C�U���4�
�<�
�$�,�$���˹��^9��V�����'�6�o�%�8�8�ǿ�&����Q��Z����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�m�3�:�j�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�e����N���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���l�3�8�m�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&����9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��@���!�0�u�u�w�}�W���YӇ��@��T��*���&�l�3�8�o�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�n�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�;�(�������V��B1�Mӊ�d�i�u����8���Hù��T9��Q��A���%�n�u�u�1��2�������l��h�� ��m�
�g�i�w�;�(�������V��X1�����3�
�a�l�'�}����	����@��A]��M��e�e�|�_�w�}�$���>����lW��C�����
� �d�b��l�K�������
]ǻN��&������!�`��(���H����CV�
N��Hԥ�l��2�4�$�8�E���&����	��R��K���|�_�u�u���;���6����9��Q��G���%�u�h�_�w�}�W�������lQ��h����u�3�
���	����O�ԓ�F9��[��E��u�u�d�|�2�.�W���Y�����Y��*���8��&�4�2���������l��h_�G�ߊu�u�����8���Aù��U��Y�����h�}�h�%�n�����
����l��D��U���0�&�k�x�~�W�W���*����v%��B��E���3�
�g�l�'�}�J�ԜY���F��G1��*��
�g�"�0�w�;�(���<����G9��h\�� ��b�
�e�e�w�}�F�������9F�N��U���;�1�
�0�:���������G��h��*���
�m�m�_�w�}�$���,����|��^��*���d�e�
�f�k�}�W���Y����`9��b"�����
�e�3�
�o��Fϩ�����V
��Z�����
�l�
�g�g�}�W��PӃ��VFǻN��U���
�d��%�#��(߁�����l�N��*����g��!�e��(���H����CW�
N��'���9�
�e�3��l�N���B��� ��O#��!ػ� �
�e�f�1��F���	���l�N��Uʳ�
���g��)�E߁�&����Q��G_�����}�0�
�8�o�4�(���H����CT�N��R��u�9�0�_�w�}�W���&�ד�]��D1��F���
�<�n�u�w�;�(���5�Ԣ�F��1��*��
�d�i�u��8����A˹��l_��h����u��-� ��3����I����V��a1�����e�
�g�i�w�)�(�������P�������1�%��&�;��@���&����CU�N�����0�}�%�6�9�)���&���9F�������;� �
�g�4�(���&����U��W�����h�&�1�9�0�>�����ι�@��R
��*��� �!�m�
�"�l�Nށ�J���F��P ��]���6�;�!�9�f��^��Y����`9��b"�����
�e�<�
�'�$��������U��N�U���u�u�u�'�#�o����ʹ��@��V�����e�`�%�u�?�3�_���&����l��Q��E���%�}�|�h�p�z�W������F�N�����%�<�
� �f�k�(��s���U5��z;��G���!�g�
�;�1�	��������l��S��U���u�u�'�!�e�4��������P��h��M���%�u�=�;��8�(���K����F9�� 1��]���h�r�r�u�;�8�}���Y���@��C�����
�b�
�f�]�}�W���������C1��D���
�a�g�%�w�`�}���Y���U5��z;��G���!�b�3�
�c�m�������@��C��*���3�
�a�c�'�u�^��^���V
��d��U���u�3�
�����������P��=N��U���-� ��;�"��(���H����CW�
N��'���9�
�d�3��i�O���B��� ��O#��!ػ� �
�
�;�2�-�!�������^��N�U���
�:�<�
�2�)�ǫ�
����WN��e�����
� �d�b��n�W�������V��G1�����9�d�
���t�L���YӀ��K+��c\�� ���
�;�3��'����O����Z�=N��U���u�0�
�
���Cށ�����R��Q��F���%�u�=�;��8�(���K����U��[�����|�h�r�r�w�1��ԜY���F��[1�����
� �d�a��n�}���Y����~3��N!��*���!�%�,�d�����O����[��d1�� ��� �
�f�d�%�:�F��B��� ��O#��!���!��9�<�;��C�������9��R�����:�&�
�#�e�n�6���8��ƹF��d1�� ����!��9�>�1�(���H����P��G^��Hʳ�
����#�l�(ށ�����^��N�������,� ��(���� ����9��hY�*��i�u�%�6�9�)���&����p"��dךU���x�2�%�3�g�;�Fށ�����l��T�����;�%�:�0�$�}�Z���YӁ��l ��h��D���
�d�
�%�4���������PF��G�����4�
�0�u�'�.��������l��h��*���4�
�<�
�$�,�$���˹��^9��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<��������]��[����h�4�
�<��.����&����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�m�3�8�`�t�^Ϫ���ƹF�N��U���'�
�
�
��l����HŹ��l��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�2�'�;�G���H¹��lQ��h�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F�	��*���
�
�d�3��l�(���
����Z�P�����3�d�
� �`�k��������R��C��*���n�u�u�2�'�;�G���H¹��lQ��h����i�u�9����4�������_��h^�����b�d�_�u�w�p�W���&����U9��h��C���4�
�0�4�$�:�W�������K��N�����3�e�3�d��(�A�������l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�d�
�&��n�W���
����@��d:�����3�8�d�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�a�3�8�f�t��������]��[����h�4�
�<��.����&����l ��h_�\���!�0�u�u�w�}�W���YӁ��l ��h��G���
�l�
�%�4�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�P�����3�d�
� �a�d�������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}�����֓�lW��Q��Lӊ�%�&�4�!�k�}����&ù��T��B1�L���
�!�'�
�'�.��������F�P�����3�d�
� �a�d��������C��R
�����`�i�u�
��<��������lV��Y1���ߊu�u�'�
���(�������
9��h>�����&�m�0�e�k�}�(؁�����V9��^ ����u�u�2�%�1�m���&����
_��Y1��9���;�
�
�
�w�`����>����l��h�����_�u�u�'���(���K����_��^ ��9���;�0�l�0�g�a�W���&����V9��1��*���n�u�u�2�'�;�G���H����lP��h��%���4�2�
�
��}�JϮ�L����T��h_�����2�_�u�u�%��(߁�&�ԓ�F9��1��*���!��
�
��}�JϽ�&����q'��X�� ���l�0�e�'�0�l�F��Y����A��h^��*���3�
�l�
�9��(���DӔ��lQ��d��Uʲ�%�3�e�3�f����@����W2��R������'�8�!�%��(ށ�����l�N�����e�3�d�
�"�k�N���&����G9��S��*ӊ�<�;�9�
��������ƹF�N�����e�3�f�3��i�(����ƭ�@�������{�x�_�u�w�/�(���&����U��Z�����
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����U�P�����3�d�
� �a�d�������R��^	������
�!�`�1�0�F���Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�}�'�>��������lW������6�0�
��$�l�(���&���R��Y��]���6�;�!�9�0�>�G������lV��h_�����l�
�%�1�9�t�^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����S��D��A���|�!�0�u�w�}�W���Y����A��h^��*ي� �c�a�4��8�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F�	��*���
�
�
� �a�i�������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}�����֓�lU��B1�A���
�!�'�u�j�:����I����l ��Z�����!�'�
�%�$�<�������F��G1��E���f�3�
�a��3�0���
�ғ�lV�
N��B���<�&�0�g�>����Y����A��h^��*ي� �c�a�<��<����&����[��hY�����
�
�
�;�$�:�}���Y����U9��Q1�����a�
�;��>�.�C���K���C9��p�����a�<�
�<�l�}�WϹ�	����l ��h��C���<�
�4�;���(���DӖ��l!��Y��*ߊ�;�&�2�_�w�}����&ù�� 9��hX�*����<�&�a�2�i�K���&Ĺ��Z��R1�����<�n�u�u�0�-�����Փ�F9��1��*���;�
�
�
�w�`����>����l��h�����_�u�u�'���(���&����R��Y1�����a�0�c�i�w��(�������9��h��N���u�2�%�3�g�;�D���&����Z��V��*ފ�
�u�h�%�`������ߓ�]9��PUךU���'�
�
�
�����M����~��V�����9�d�
�
�w�`����4����_%��C��*���
�;�&�2�]�}�W���&����U9��Q��Aފ�;��;�4��3����H����F���*��� �9�:�!�8��(ށ�����l�N�����e�3�f�3��i�(���4����_%��C��*���0�g�i�u����������A	��R1�����<�n�u�u�0�-�����Փ�F9��1��*��� �9�:�!�8��E���J���C9��z�����;�'�9�0�d�4�(���B�����h��*���
� �c�a�>���������A	��\��*���h�%�a��9�<�4�������lR��Y1���ߊu�u�'�
���(܁�����l��z�����;�'�9�d���W��	�ғ�R��[-�����
�
�
�;�$�:�}���Y����U9��Q1�����a�
�;��9�<�4�������9��N�U���
�4� �9�8�)����&Ź��l��d��Uʲ�%�3�e�3�d�;�(��&����R��[-�����
�g�0�b�k�}�(ہ�����p	��E�����<�
�<�n�w�}�����֓�lU��B1�A���
��g�0�g�a�W�������G��h:�����4�0��
�%�����N����F�P�����3�f�3�
�c�����&����F���D���%�!�
�
��3����s���T��Q1�����3�
�a�
�9��(݁�&��� ��O/�����
�d�d�'�0�l�@��Y����A��h^��*ي� �c�a�<���E���J���U5��d;��:����7�'�6��e�F�������
]ǻN�����
�
�
�
�"�k�C���&����V9��R1�I���
�
�4�2���(���
����F�P�����3�f�3�
�c���������l��R������;�0�0�d�4�(���B�����h��*���
� �c�a�>�����&Ĺ��F���*���2�
�
�
�9�.��ԜY�ƫ�C9��1��F���
�a�
�;��3�������F��1�����0�`�<�
�>�f�W�������lV��h]�� ��a�<�
�4�0��(���Y����lS��V ��*���
�;�&�2�]�}�W���&����U9��Q��Aފ�;��;�0�`�8�B��Y����a��R1��B���
�<�n�u�w�:����I����l ��Z�����4�2�
�
��}�JϮ�L����T��hV�����2�_�u�u�%��(߁�&����lP��h��'���0�b�0�b�k�}�(ځ�����V9��^ ����u�u�2�%�1�m��������9��h=��D���e�i�u�
��<��������lV��Y1���ߊu�u�'�
���(܁�����l��d>��*���u�h�%�d��8��������9��h��N���u�2�%�3�g�;�D���&����Z��R��*���h�%�l��0�<����H����@��=d��U���u�'�
� �`�h����
������T��[���_�u�u�'��(�@�������@��h����%�:�0�&�6�����
����g9��1����u�%�6�y�6�����
����g9��1����u�%�&�2�4�8�(���
�ߓ�@��N��*���
�&�$���)�C���������h=�����
�
�
�0�3�/��������l�������6�0�
��$�o�(���&���R��^	������
�!�`�1�0�E������T9��R��!���d�
�&�
�a�}��������B9��h��@���8�d�y�2�'�;�G���J����R��V�����u�%�&�2�4�8�(���
����U��W����<�
�&�$����������J��G1�����0�
��&�f�����L�ƭ�l��h�����
�!�l�3�:�l�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y����\�V�����
�:�<�
�w�}����P�ƣ�N��h�����:�<�
�u�w�-��������`2��CV�����|�:�u�4��2��������F�V�����&�$��
�#�����PӉ����T�����2�6�d�h�6�����
����g9��Z�����f�u�'�}�'�>��������lW������6�0�
��$�o�(���&���\�V�����
�:�<�
�w�}��������B9��h��@���8�g�|�:�w�u��������\��h_��U���&�2�6�0��	���&����R�V ��]´�
�:�&�
�!��W���&ʹ��T��D1��G���4�
�0�1�1��N݁�K�ƣ�N��h�����:�<�
�u�w�/�(���&����U��Z�����;�|�|�:�w�u��������EW��S��*ӊ�<�;�9�
����������U��\��G���;�u�4�
�8�.�(�������F��h��*���$��
�!�a�;���P�ƣ�N��G1�����9�d�e�h�'�d�$�������lT��R�����
� �g�g�'�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���'�}�4�
�8�.�(���&���C9��d�����0�g�'�4��8����&����CT�V ��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�`�t����Q����\��h��*���u�
�
�<�9�1�(���&����l��S1��*��
�g�u�;�w�<�(���
����T��N�����<�
�&�$����������O�X��]���6�;�!�9�f�m�JϮ�@����]��h��*���1�'�4�
�"�o�E���PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����d�|�|�u�?�3�}���Y���F�P�����g�
�0�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����A��B1�@���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���'�
� �b�b�2����Y����T��E�����x�_�u�u�%����L����\��V�����'�6�o�%�8�8�Ǯ�@����]��h��*���1�'�4�
�"�o�E���UӇ��@��T��*���&�d�
�&��q��������V��c1��Dߊ�&�
�a�u�'�.��������l��1����y�4�
�<��.����&����U��B�����2�6�0�
��.�B������R��^	������
�!�d�1�0�F������T9��R��!���d�
�&�
�`�}��������B9��h��G���8�g�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�b�}����	����@��X	��*���u�%�&�2�4�8�(���
�ԓ�@��N��U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ԓ�@��G�����:�}�4�
�8�.�(���&���C9��d�����0�g�'�4��8����&����CT���U´�
�:�&�
�8�4�(���Y����Z��D��&���!�`�3�8�f�t�^������F�N��U���2�%�3�
�e��������R��X ��*���
�n�u�u�w�}�������R��X ��*���<�
�u�u�'�.��������l��1����u�'�}�%�4�3��������[��G1�����0�
��&�f�����I�ƣ�N��CF�����;�!�9�d�g�`����*����_��h\�����'�4�
� �e�o����Y������T�����2�6�d�h�6�����
����g9��V�����b�|�|�!�2�}�W���Y���F��E�� ��`�:�6�1�w�`��������_��UךU���u�u�9�0�]�}�W���Y���T��Q��Gߊ�%�:�0�i�w��U�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�P�����g�
�e�4�$�:�W�������K��N�����3�
�g�
�g�<����&����\��E�����
�d��%�#��(ށ�����F��P1�L���0�
�e�y�%�:�O��Y����~3�� ����
�
�0�
�`�l�W���
����@��d:�����3�8�l�u��%�"���6����F
��G��C���'�2�d�c�{�<�(���&����l5��D�*���
�a�u�%�$�:����&����GT��Q��G���2�%�3�e�1�n����Mǹ��l��B��L���%�&�2�6�2��#���K����lW�V�����&�$��
�#�����UӇ��@��T��*���&�d�
�&��m�W���
����@��d:�����3�8�d�y�6�����
����g9��\�����d�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��G܊�&�
�`�|�#�8�W���Y���F�	��*���b�`�%�u�j�/���@���F�N�����}�4�
�:�$�����&���R��^	������
�!�m�1�0�F���Y����l�N��U���u�2�%�3��o�(��E�ƾ�T9��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����R����ߊu�u�u�u�w�}��������l��S�����
�
�
�
�"�k�C���&����A��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�:����&����CV�
N��*����,� �
�"�)����O�ד�V�� X����u�u�u�9�>�}�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����֓�@��N��U´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�e�t�^Ϫ���ƹF�N��U���'�
� �b�b�-�W������R��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�2�'�;�(��&���F��_�����&�0�d�<��4�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�~�)����Y���F�N����� �b�`�%�w�`����4����])��h\��D���2�d�e�n�w�}�W�������9F�N��U���u�'�
� �`�h����D�Ĕ�k>��o6��-���������/���!����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʲ�%�3�
�g��l�����Ƽ�\��D@��X���u�2�%�3��o�(�������]9��X��U���6�&�}�
�f�����&����Z��^	���
�;� �&�2�o��������V�� ]����b�l�u��/��#�������G��N1��D���2�d�`�y�6�����
����g9��^�����y�4�
�<��.����&����l ��h_�U���-� ��;�"��(ށ�����R�V�����&�$��
�#�k����K����C9��P1������&�g�3�:�l�W���
����@��d:��ߊ�&�
�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
����U��Y����<�
�&�$����������OǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����Г�@��G�����u�u�u�u�w�}�WϹ�	����T��G_��Hʳ�
���g��)�@�������Q��=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�Fׁ�
����O��_�����u�u�u�u�w�/�(���N�ӓ�F���*��n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����W��D��E���!�0�u�u�w�}�W���YӁ��l �� \�����h�3�
���$��������_��h_�����b�g�_�u�w�}�W��������T�����2�6�d�h�6�����
����g9��^�����|�:�u�4��2��������F�V�����&�$��
�#�h����H����AF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�d�|�u�?�3�}���Y���F�P�����g�
�d�i�w�8�(��B���F������}�%�6�;�#�1����H����C9��P1������&�`�3�:�i�^Ϫ���ƹF�N��U���'�
� �b�b�-�W��	����z��C��*؊�;�&�2�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C\�����|�u�=�;�]�}�W���Y���T��Q��Gߊ�d�i�u�
�f�����&����Z��^	�U���u�u�0�&�w�}�W���Y�����h��B���%�u�h�w���/���!����k>��o6��-������w�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƫ�C9��hY�*���4�&�2�u�%�>���T���F��G1��*��
�0�4�&�0�����CӖ��P�������6�0�
��$�l����I�ƭ�l�������6�0�
��$�e����N�ƭ�l��h�����
�!�
�&��q��������V��c1��Dފ�&�
�f�u����������9��V
�����3�
�l�
�e�}��������B9��h��D���8�g�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
����U��X����<�
�&�$����������J��E��*ڊ�
�
� �c�c�<�(����ƭ�l��h�����
�!�e�3�:�l�[Ͽ�&����P��h=����
�&�
�b�w�-��������`2��C_�����d�y�4�
�>�����*����_��D��M�ߊu�u�0�<�]�}�W���Y���N��h�����:�<�
�u�w�-��������`2��C_�����|�:�u�:��<�(���
����T��N�����0�|�:�u�6�����&����P9��
N��*���
�&�$���)�(���&����AF��G1�����9�2�6�d�j�<�(���&����l5��D�����m�u�'�}�'�>��������lW������6�0�
��$�l�(���&���\�V�����
�:�<�
�w�}��������B9��h��D���8�g�|�:�w�<�(���
����T��N�����<�
�&�$����������O��EN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�l�w�/�_�������l
��^��U���%�&�2�6�2��#���H˹��^9��N��U���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��i�W���Y�έ�l��D��ۊ�u�u�
�
�>�3����&����R��R�����l�
�g�u�%�u��������\��h^��U���
�
�
�
��(�A�������]�N��U���%�6�;�!�;�l�G��	�ߓ�Z��[��*؊�0�1�'�4��(�E���	����]�V�����
�:�<�
�w�}��������B9��h��C���8�d�|�u�%�u��������_��N������2�4�&�2�o����&����l ��W�����4�1�}�%�4�3��������[��G1�����0�
��&�f�����O����AF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�m�|�u�?�3�}���Y���F�P�����g�
�0�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����A��B1�L���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���'�
� �b�n�2����Y����T��E�����x�_�u�u�%����@����\��V�����'�6�o�%�8�8�Ǯ�@����]��h��*���1�'�4�
�"�o�E���UӇ��@��T��*���&�d�
�&��q��������V��c1��Dߊ�&�
�a�u�'�.��������l��1����y�4�
�<��.����&����U��B�����2�6�0�
��.�B������R��^	������
�!�d�1�0�F������T9��R��!���g�
�&�
�f�W�W�������F�N�����}�4�
�:�$�����&���R��^	������
�!�e�1�0�N����έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���:�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������C9��Y�����6�d�h�4��4�(�������@��Q��A���'�}�%�6�9�)���������D�����
��&�d��.�(��P�Ƹ�V�N��U���u�u�2�%�1��Eց�	����Z�V�����
�#�
�n�w�}�W�������N�V�����
�:�<�
�w�}��������B9��h��G���8�g�|�:�w�3����	����@��A_��U���
�
�<�;�;��(݁�����V��Q��L؊�g�|�4�1��-��������Z��S�����2�6�0�
��.�Fځ�
����O����ߊu�u�u�u�w�}��������l	��X
��I���%�6�;�!�;�o�G�ԜY���F��D��U���u�u�u�u�0�-����Kʹ��P	��R��W���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������
9�������%�:�0�&�w�p�W�������F9��1��*���<�;�%�:�w�}����
�ξ�T9��B�����l�y�3�
���E������� 9��P1�E���4�
�<�
�$�,�$����֓�@��N��*����,� �
�"�)����H����A��Y�Yʴ�
�<�
�&�&��(���L����lW����;����!�d�
�"�l�Oց�H�ƭ�l��h�����
�!�c�3�:�o�[Ͽ�&����P��h=�����3�8�d�u�'�.��������l��h��*���4�
�<�
�$�,�$����ד�@��B�����2�6�0�
��.�E݁�
����l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���KŹ��^9��G�����_�u�u�u�w�}�W���&����_��N�U������!�f����Aʹ��l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�l����H���G��d��U���u�u�u�2�'�;�(��&���F��h��9��� �
� �!�'�$�F݁�&����Q��d��U���u�0�&�3��u��������\��h_��U���&�2�6�0��	���&����
O��EN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�a�w�/�_�������l
��^��U���%�&�2�6�2��#���K����^9��G�����u�u�u�u�w�}�WϹ�	����T��G^��Hʧ�2�b�b�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C[�����|�u�=�;�]�}�W���Y���T��Q��Gӊ�e�i�u�0��j�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�~�)����Y���F�N����� �b�l�%�w�`����4����])��h\��F���2�d�e�n�w�}�W�������9F�N��U���u�'�
� �`�d����D�Ĕ�k>��o6��-���������/���!����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʲ�%�3�
�g��l�����Ƽ�\��D@��X���u�2�%�3��o�(�������]9��X��U���6�&�}�
�f�����&����Z��^	���
�;� �&�2�i��������V��W����<�
�&�$����������F��h��9��� �
� �!�'�$�Fځ�&����Q��N��*���
�&�$���)�B������� ��O#��!ػ� �
�
�
�2��O��Y����Z��D��&���!�c�3�8�e�q�����֓�lU��B1�A���
�0� �;�o�}��������B9��h��*���
�y�4�
�>�����*����9��Z1�U���&�2�6�0��	���&����V�V�����&�$��
�#�o����K��ƹF��R	�����u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�:����&����CW�
N��*����g��!�`�l����H����9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����M����[��=N��U���u�u�u�'��(�@���	�����h��*���
� �c�a�6���������F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!�f�;���P�Ƹ�V�N��U���u�u�2�%�1��Eց�H���U5��z;�����
� �!�%�.�l�(ށ�����Q��N��U���0�&�3�}��-��������Z��S�����2�6�0�
��.�F߁�
����	�������!�9�2�6�f�`��������V��c1��G؊�&�
�d�|�w�5��ԜY���F�N�����
�g�
�d�k�}����I��ƹF�N�����u�}�%�6�9�)���������D�����
��&�`�1�0�C�������9F�N��U���u�'�
� �`�d����DӖ��9��G��*���
�;�&�2�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��G1��*��
�d�i�u��l�>�������9��h��N���u�u�u�0�$�}�W���Y���F��E�� ��l�%�u�h�u��/���!����k>��o6��-�������u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���T��Q��Fي�0�4�&�2�w�/����W���F�P�����f�
�0�4�$�:�(�������A	��D�����y�4�
�<��.����&����U��B�����2�6�0�
��.�B������R��^	������
�!�
�$��^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�4�
�8�.�(�������F��h��*���$��
�!��.�(�������C9��Y�����6�d�h�4��4�(�������@��Q��A���'�}�%�6�9�)���������D�����
��&�c�1�0�B���PӒ��]FǻN��U���u�u�'�
�"�j�D���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʲ�%�3�
�f��8�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�2�'�;�(��&���F��_�����&�0�a�<��4�L���YӁ��l �� ]�����h�%�d�
�9�(����L����@��=d��U���u�'�
� �`�j����
������T��[���_�u�u�'��(�@�������@��h����%�:�0�&�6�����	����l��F1��*���
�&�
�y�6�����
����g9��1����u�%�&�2�4�8�(���
�Г�@��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}����Q����\��h�����u�u�%�&�0�>����-����l ��hX�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t��������]��[����h�4�
�<��.����&����U��G��\ʡ�0�u�u�u�w�}�W�������F9�� 1��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������l��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�ƫ�C9��hY�*��i�u�0�
�o�f�W�������F9�� 1��U��%�d�
�;�"�.��������T]ǑN��X���'�
� �b�d�-�W�������A	��D�X�ߊu�u�'�
�"�j�D���&����T��E��Oʥ�:�0�&�'�0�j�D�������
J��G1�����0�
��&�o�;���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�*���
�f�u�%�$�:����&����GT��Q��G���4�
�<�
�$�,�$����ӓ�@��B�����d�y�3�
������&����Z��h_��D���2�d�a�y�6�����
����g9��^�����y�3�
������&¹��T9�� \������� ��m�E�������OǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ӓ�@��G�����u�u�u�u�w�}�WϹ�	����R��G^��Hʧ�2�m�a�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C\�����g�|�u�=�9�W�W���Y���F��G1��*��
�e�i�u���;���6����9��E��D���n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����R��D��F���!�0�u�u�w�}�W���YӁ��l �� Z�����h�3�
������&¹��T9�� \�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���I����l_����ߊu�u�u�u�w�}��������l��S��&��� ���!��1����&�ѓ�l��h_�E�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ߓ�@��G�����_�u�u�u�w�}�W���&����U��N�U���
�m�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y����A��B1�F���u�h�'�2�`�n�}���Y���V
��d��U���u�u�u�2�'�;�(��&���F��o6��-���������/���!����k>�=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�'�
�"�j�D���Y����T��E�����x�_�u�u�%����J����R��P �����o�%�:�0�$�-�A�������V��R1�����<�y�4�
�>�����*����9��Z1�U���&�2�6�0��	��������F��h��*���$��
�!�c�;���UӇ��@��T��*���&�g�
�&��m�W���
����@��d:�����3�8�g�y�1���������@��X��9���g�
�0�
�`�e�W���
����@��d:�����3�8�l�_�w�}����s���F�^��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�c�t����Y���F�N��U���
� �b�f�'�}�JϿ�&����G9��\��3ߑ�a�e�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���T��Q��Aي�d�i�u�
��<��������lU��Y1���ߊu�u�u�u�;�4�W�������]��[����h�4�
�<��.����&����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��m�W���Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����U��]��D��u��;�1��8��������t*��h\�����d�g�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y����A��B1�F���u�h�4�
�8�.�(���K�Պ� %��UךU���u�u�9�0�]�}�W���Y���T��Q��Aي�d�i�u����/���!����k>��o6��-������n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӁ��l �� Z�����&�<�;�%�8�8����T�����h��B���%�
�&�<�9�-����Y����V��E��B��u�0�
�m�{�<�(���&����l5��D�����b�u�%�&�0�>����-����l ��hV����<�
�&�$���������� J��G1�����0�
��&�e�����I�ƪ�l��{:�� ��� �!�%�,�f��(���&����F��h��*���$��
�!�g�;���Y����`3��x��&���'�6�
�m�f�/���N����`9��{+��:���m�
�
�0��e�C�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����I����[��=N��U���u�u�u�'��(�@���	��� ��d+��6���!�m�
�
�2��O��s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�a�3�:�l�^������F�N��U���2�%�3�
�c��G��Y����`3��x��&���'�6�
�m�f�/���N��ƹF�N�����u�}�%�6�9�)���������D�����
��&�d��.�(���Y����l�N��U���u�2�%�3��i�(��E�ƪ�l��{:�� ��� �!�%�,�f��(���&����l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�2�%�1��Cׁ�I���A�� V����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���A����lQ����ߊu�u�u�u�w�}��������l��S�����m�n�u�u�w�}����Y���F�N��U���
� �b�m�'�}�J���!����k>��o6��-���������/���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����
�a�
�d�6�.��������@H�d��Uʲ�%�3�
�a��l��������\������}�
�
�4�6�8�����Փ�]9��PB�����2�6�0�
��.�O������R��^	������
�!�
�$��[Ͽ�&����P��h=����
�&�
�f�w�-��������`2��C\�����g�y�3�
�8�8����&����\��{��Gۊ�0�
�b�a�w�-��������`2��C_�����l�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��Dފ�&�
�f�|�#�8�W���Y���F�	��*���b�m�%�u�j�-�A�������V��R1�����<�n�u�u�w�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���:�u�4�
�8�.�(�������F��h��*���$��
�!�f�;���PӉ����T�����2�6�d�h�6�����
����g9��^�����|�|�!�0�w�}�W���Y�����h��B���%�u�h�3��2��������]��d)����
�0�
�b�c�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:��Ҋ�&�
�|�u�?�3�}���Y���F�P�����a�
�d�i�w�-��������9��v/��4��u�u�u�u�2�.�W���Y���F�	��*���b�m�%�u�j��/���!����k>��o6��-���������}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��G1��*���
�e�4�&�0�}����
���l�N�����
�`�
�e�6�.���������T��]���&�2�6�0��	��������F��h��*���$��
�!�f�;���UӔ��lQ��N��*����,� �
�"�)����Hǹ��A��Y�Yʴ�
�<�
�&�&��(���I����l_�Q=��0���� �
�c�e�/���O��ƹF��R	�����u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�:����&����CV�
N��*����� �
�a�o����H����9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����P�Ƹ�V�N��U���u�u�2�%�1��B܁�I���U5��z;�����
� �!�%�.�l�(ށ�����P��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�2�'�;�(��&���F��P1�B�ߊu�u�u�u�;�8�}���Y���F�P�����`�
�e�i�w��/���!����k>��o6��-��������f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӁ��l �� [�����h�3�
�:�2�)��������`!��^1�*���
�b�a�_�w�}�Z�������lQ��h����2�u�'�6�$�s�Z�ԜY�ƫ�C9��hY�*���4�&�2�
�%�>�MϮ�������D�����
��&�l�1�0�O���	����l��F1��*���d�3�8�g�{�/���N�ƪ�l��{:�� ��� �!�%�,�f��(���&����F��h��*���$��
�!�g�;���Y����v*��c!��*���g�'�2�d�a�t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�d�1�0�E���Y����l�N��U���u�2�%�3��h�(��E�ƪ�l5��r-�� ���c�g�'�2�f�k�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�~�}����s���F�N�����3�
�`�
�g�a�W�������J)��h#�����,�d�
�
�2��@��s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��Uʲ�%�3�
�`��m�K�������]ǻN��U���9�0�_�u�w�}�W���Y����U��Y��E��u������/���!����k>��o6��-����n�u�u�w�}�������F�R �����0�&�_�u�w�:����&����CW�
N��*���0�!�'�
�>�>��������l��h_�M�ߊu�u�:�
��d����Jƹ��Z�G1��؊�
� �m�d�'�u�D��Hӂ��]��G�U���9�6��g��(�F��&���F��a��*���3�
�e�d�'�u�GϺ�����U�=N��U���
�
�d�3��m�B���Y����l0��1�*���d�d�
�d�e�}�W�������V�=N��U���
�
�g�3��o�C���Y����l0��1�*���d�l�
�d�d�}��������l�N�����g�
� �d�g��F��Y����_T��1��*��d�%�}�f�z�l��������l�N�����3�
�g�
�c�a�W����ԓ�l ��\�����e�1�"�!�w�n�L���YӖ��V��1��*���d�g�
�f�k�}�W���Y����C9��Y����
�u�=�;��0�(�������Q��F�U���d�|�0�&�w�}�W���Yӊ��l0��1��*��`�%�n�u�w�-�G��&¹��l ��Z�*��i�u�u�u�w�}��������_��h^�����}�8�
�a�1��D���	����[�I�����u�u�u�u�w�1����K����lW��1��N���u�%�e�e���(���@�Փ� F�d��U���u�4�
�:�$�����Iӑ��]F��Z�� ��b�%�}�|�j�z�P������F�N������d�
� �o�h���Y����lV��T�����
�u�h�6��2��������A��_��%���&�6�d�'�0�l�O��s���K��h^�����;�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�e��)�����֓�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!�o�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���F��R ��U���u�u�u�u�'�m�6�������lV��G1����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����8����]��h^�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN������!�:�&�2�l�K�������V9��E������4�0���/�(݁�����
W��=N��U���%�e��!�8�.��������WF��D��U���6�&�{�x�]�}�W���&����\��R1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K˹��^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h\�\���=�;�_�u�w�}�W���Y����r��X �����4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��v�����0�d�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
��>����&����[��[1�����0�8��&�6�8�4�������l��h_�G�ߠu�u�x�u����������9��h��U���<�;�%�:�2�.�W��Y����lV��T�����
�
�%�#�3�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����g�|�|�!�2�}�W���Y���F��h^�����;�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8����Y���F�N��*ڊ�6�<�;�
���������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����8����]��h]��Hʶ�
�:�0�!�%���������]��[1��D���2�d�e�n�]�}�W��	�֓�P��Y��*ي�%�#�1�4�$�:�W�������K��N������!�:�&�2�n��������@��h����%�:�0�&�6�����	����l��F1��*���m�3�8�g�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��j�^������F�N��U���%�e��!�8�.��������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�e��)�����Փ�C9��SN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���C9��v�����0�a�i�u�;�3��������R��S�����:�
�
�
�2��O��s���K�G1��4���:�&�0�a�6�����
������T��[���_�u�u�
��>����&����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�����N���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�O�������O��_�����u�u�u�u�w��(�������V9��V�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����\��R1�����9�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=N��U���
�6�<�;���W������W��R��6���4�0��;�%�1��������W��=d��U���u�
�
�6�>�3�(���&����_��D��ʥ�:�0�&�u�z�}�WϮ�I����Z	��h��*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ޓ�@�� GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӖ��l'��^��*���
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����h/�����
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�%�g�����
����Z�T�����!�'�
�4�4�9��������@9��E��D��n�_�u�u�z�-�G�������l��h�����4�&�2�u�%�>���T���F��1�����&�0�c�4��1�(�������A	��N�����&�4�
�0�w�-��������`2��C\�����g�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��GҊ�&�
�b�|�w�5��ԜY���F�N��E���!�:�&�0�a�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�e��!�:�$�8�A���&����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���&ù��G��D1��B��u�9�;�1��8����
����W%��C��*���
�0�
�m�`�W�W���T�Ƽ�9��C�����b�4�
�9�w�.����	����@�CךU���
�
�6�<�9��(؁�	����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�g�
�&��j�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�m�1�0�E���PӒ��]FǻN��U���u�u�
�
�4�4����&Ĺ��l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u����������9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��h^�����;�
�
�u�j�>�(�������^9��D�����;�'�9�&�a�/���J��ƓF�C��*ڊ�6�<�;�
������Ӈ��Z��G�����u�x�u�u�'�m�6�������l^��G1�����&�2�
�'�4�g��������C9��N��*���
�&�$���)�O�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����Q�N�����u�u�u�u�w�}����8����]��hV�����1�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W���	�֓�P��Y��*Ҋ�%�#�1�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%�e��!�8�.���E�Ư�l��R1�����4�6�1�1�8�)����&Ĺ��T9��Y����u�x�%�e��)�����ߓ�C9��SN�����u�'�6�&�y�p�}���Y����r��X �����4�
�9�
�$�4��������C��R�����0�u�%�&�0�>����-����9��Z1�\���u�7�2�;�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�]�}�W���Y���C9��v�����0�l�4�
�;�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�G1��4���:�&�0�l�6�����DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���I����C	��C��*ڊ�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�e��)����
����l��A�����<�
�&�<�9�-����Y����V��G1�*���%�<�!�
�������Ƽ�V��R�����
�
�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��Dڊ�0�%�<�!���(��������YNךU���u�u�u�u��m�$�������l��h�����<�
�<�u�j�-�F߁�����]��R1�����9�n�u�u�w�}����Y���F�N��U���e��!�:�9�.��������W9��h��U��%�d�
�0�'�4����&ù��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��G�������G��h^�����2�4�&�2�w�/����W���F�G1�*���%�<�!�
����������Z��G��U���'�6�&�}��m�$�������l��N��Dڊ�0�%�<�!���(����Ƽ�V��R�����
�
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������1�����;�&�0�e�6�����Y����l�N��U���u�%�d�
�2�-����&����Z��^	��Hʥ�d�
�0�%�>�)�(���B���F����ߊu�u�u�u�w�}�(���*����Z��h��*���&�2�i�u��m�$�������l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��F���	����V9��V�����;�&�2�4�$�:�W�������K��N����
�;� �&�2�m��������l��h�����%�:�u�u�%�>����&�ד�]��D1��E���
�9�y�%�f�����
����l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(���0����@9��1��*���|�u�=�;�]�}�W���Y���C9��h'�� ���0�e�4�
�;��������C9��h'�� ���0�e�4�
�;�f�W���Y����_��=N��U���u�u�u�
�f�����&����R��[
�����2�i�u�
�f�����&����R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(���0����@9��1��*���u�&�<�;�'�2����Y��ƹF��h_��<���!�
�
�
�9�.����
����C��T�����&�}�
�d��-����&����lW��~ �����
�
�'�2�w��F���	����V9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��F���	����V9��V�����u�=�;�_�w�}�W���Y�Ƽ�W��Y�����e�<�
�<�w�`���&����G��h^�U���u�u�0�&�w�}�W���Y�����1�����
�
�
�;�$�:�K���&�ד�]��D1��E���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�H¹��C��h��*���#�1�<�
�>�}����Ӗ��P��N����u�
�d��'�)�(���&����_��Y1�����&�2�
�'�4�g��������lW��~ �����
�
�%�#�3�}�(���0����@9��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	����z��C��*ۊ�%�#�1�|�#�8�W���Y���F���D���%�!�
�
��-��������TF���D���%�!�
�
��-����s���F�R��U���u�u�u�u�w�-�Fށ�����l��h�����<�
�<�u�j�-�Fށ�����l��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	����z��C��*ۊ�;�&�2�4�$�:�W�������K��N����
�;� �&�2�l��������@��h����%�:�0�&�'�l�(�������lW�G1�*��� �&�0�d�'�8�[Ϯ�H¹��C��h��*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�H¹��C��h��*���#�1�|�!�2�}�W���Y���F��h_��<���!�
�
�
�9�.���Y����l/��B����_�u�u�u�w�1��ԜY���F�N��Dۊ�;� �&�0�f�4�(���Y����lW��~ �����
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�W��Y�����g�4�
�9��3��������]F��X�����x�u�u�%�f�����
����l��A�����<�
�&�<�9�-����Y����V��G1�*��� �&�0�g�6����	����z��C��*؊�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��h'�� ���0�g�4�
�;�t�W������F�N��Uʥ�d�
�;� �$�8�E���&����Z��^	��Hʥ�d�
�;� �$�8�E���&����9F�N��U���0�_�u�u�w�}�W���&�ד�]��D1��G���
�9�
�;�$�:�K���&�ד�]��D1��G���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��h'�� ���0�g�<�
�>�}����Ӗ��P��N����u�
�d��'�)�(���&����Z��D�����:�u�u�'�4�.�_���H����F��R1�U���d��%�!���(����Ƽ�W��Y�����g�4�
�9�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�W��Y�����g�4�
�9�~�}����s���F�N����
�;� �&�2�o���������1�����
�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�d��%�#��(݁�����Z�G1�*��� �&�0�g�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h_��<���!�
�
�
�'�+����&����R��P �����&�{�x�_�w�}�(���0����@9��1��*���
�;�&�2�6�.���������T��]���d��%�!���(������C9��h'�� ���0�f�4�
�;�����s���Q��Yd��U���u�<�u�}�'�>��������lW���D���%�!�
�
��-����PӒ��]FǻN��U���u�u�
�d��-����&����l��h�����i�u�
�d��-����&����l��d��U���u�0�&�u�w�}�W���Y����lW��~ �����
�
�%�#�3�4�(���Y����lW��~ �����
�
�%�#�3�-���Y���F��Y
�����u�u�0�1�'�2����s���F���D���%�!�
�
��3��������]F��X�����x�u�u�%�f�����
����l��D�����2�
�'�6�m�-����
ۖ��9��G��*���y�%�d�
�9�(����J����TJ��h_��<���!�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h_��<���!�
�
�
�'�+��������9F�N��U���u�
�d��'�)�(���&����Z�
N��Dۊ�;� �&�0�d�W�W���Y�Ʃ�@�N��U���u�u�%�d��3�����Փ�]9��PN�U���d��%�!���(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C���
�;� �&�2�i��������l�������%�:�0�&�w�p�W���	����z��C��*ފ�%�#�1�<��4�(�������A	��N�����&�%�d�
�9�(����M����E
����D���%�!�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�d�
�;� �$�8�C���&����F��R ��U���u�u�u�u�'�l�(�������lR��G1�����
�<�u�h�'�l�(�������lR��G1���ߊu�u�u�u�;�8�}���Y���F�G1�*��� �&�0�a�6���������Z�G1�*��� �&�0�a�6���������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�d�
�;� �$�8�C���&����R��P �����&�{�x�_�w�}�(���0����@9��1��*���
�&�<�;�'�2�W�������@N��_�����&�0�a�u��l�>�������9��R	���
�;� �&�2�i������ƹF��R	�����u�u�u�3��<�(���
����T��N����
�;� �&�2�i�������G��d��U���u�u�u�%�f�����
����l��D��I���
�d��%�#��(��Y���F��[�����u�u�u�u�w��F���	����V9��^ �����h�%�d�
�9�(����M����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�d��'�)�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��h'�� ���0�`�4�
�;���������Z��G��U���'�6�&�}��l�>�������9��h��Yʥ�d�
�;� �$�8�B���&����C��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�d��-����&ƹ��l��G�����_�u�u�u�w�}�W���H����F��R1�����9�
�;�&�0�a�W���H����F��R1�����9�n�u�u�w�}����Y���F�N��U���d��%�!���(�������]9��PN�U���d��%�!���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�d��-����&ƹ��l�������%�:�0�&�w�p�W���	����z��C��*ߊ�;�&�2�4�$�:�(�������A	��D��*����%�!�
��q���&����G��h[�����u�
�d��'�)�(���&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�d��'�)�(���&����_����ߊu�u�u�u�w�}�(���0����@9��1��*���u�h�%�d��3��������F�N�����u�u�u�u�w�}�WϮ�H¹��C��h��*���&�2�i�u��l�>�������9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�f�����
����l��A�����<�u�&�<�9�-����
���9F���D���%�!�
�
��-��������T9��D��*���6�o�%�:�2�.���&����G��hX�����1�u�
�d��-����&Ź��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�l�(�������lP��G1�����!�0�u�u�w�}�W���YӖ��9��G��*���
�%�#�1�>�����DӖ��9��G��*���
�%�#�1�]�}�W���Y����l�N��U���u�%�d�
�9�(����O����E
��^ �����h�%�d�
�9�(����O����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�l�(�������lP��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��h'�� ���0�c�<�
�>���������PF��G�����%�d�
�;�"�.���Y����l/��B�����%�0�y�%�f�����
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�f�����
����l��A��\ʡ�0�u�u�u�w�}�W���	����z��C��*܊�;�&�2�i�w��F���	����V9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�W��Y�����c�<�
�<�w�`���&����G��hX�����_�u�u�u�w�3�W���Y����������n�_�u�u����������F������,� �
�
�2��O��s���K�G1��:��� �&�0�e�6�����
������T��[���_�u�u�
��(����&����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�����N���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�O�������O��_�����u�u�u�u�w��(���	����V9��V�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����F��R1�����9�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=N��U���
� �%�!���W������F9��1��N���u�%�f��#�(����H�����q+��7���:�!� �
�n�8�G�������]ǑN��X���
�
� �%�#��(�������WF��D��U���6�&�{�x�]�}�W���&����F��R1�*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ޓ�@�� GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӖ��l)��G��*���e�4�
�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��1�����&�0�d�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����6����G��h_�����1�4�&�2�w�/����W���F�G1��:��� �&�0�d�6�����
����l��TN����0�&�4�
�2�}��������B9��h��M���8�g�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�b�~�}����s���F�N������!� �&�2�l���������T�����2�6�d�_�w�}�W������F�N��U���%�f��!�"�.��������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����|��B����i�u�'�
�"�j�N���B���F���*���%�!�
�
��-��������]F��X�����x�u�u�%�d�����
����l��A�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�e����K��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Eׁ�
����O�C��U���u�u�u�u�w�-�D�������l��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�J����C��h��*���#�1�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʥ�f��!� �$�8�D��Y����`3��x��L���2�d�c�n�]�}�W��	�Փ�F��C��*ي�%�#�1�4�$�:�W�������K��N������!� �&�2�n��������@��h����%�:�0�&�6�����	����l��F1��*���m�3�8�g�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��j�^������F�N��U���%�f��!�"�.��������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�f��)�����Փ�C9��SN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���C9��x�� ���0�a�i�u�2��F��s���K��h]�� ���!�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�f��)�����ғ�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!�o�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���F��R ��U���u�u�u�u�'�n�8�������lR��G1����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����6����G��hZ�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN������!� �&�2�h�K������� ]ǑN��X���
�
� �%�#��(ځ�	������^	�����0�&�u�x�w�}����6����G��h[�����1�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���A����lT��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��Y��\ʡ�0�u�u�u�w�}�W���	�Փ�F��C��*ߊ�%�#�1�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����lU��B�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�f��)�������F��P1�D�ߠu�u�x�u����������9��h��U���<�;�%�:�2�.�W��Y����lU��B�����
�
�%�#�3�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����g�|�|�!�2�}�W���Y���F��h]�� ���!�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8����Y���F�N��*ي� �%�!�
���������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����6����G��hY��Hʳ�
����#�o�(ށ�����T��=N��U���%�f��!�"�.��������WF��D��U���6�&�{�x�]�}�W���&����F��R1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K˹��^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h\�\���=�;�_�u�w�}�W���Y����|��B�����4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��x�� ���0�b�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
��(����&����[��d1�� ��� �
� �!�6�)�Fׁ�&����Q��dךU���x�%�f��#�(����A����E
��V�����'�6�&�{�z�W�W���&����G��D1��M���
�9�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��Y��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����^��D��B���u�=�;�_�w�}�W���Y�Ƽ� 9��C�����m�4�
�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��1�����&�0�m�4��1�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u����������
F������
�0�8��%�8����)����A��R	��B��_�u�u�x�w��(���	����V9��V�����&�<�;�%�8�8����T�����h!�����
�
�
�%�!�9��������\������}�%�6�y�6�����
����g9��V�����b�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��M���8�g�|�|�#�8�W���Y���F���*���%�!�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���
� �%�!���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l+��B�����:�
�
�
�'�+����&����R��P �����&�{�x�_�w�}�(ہ�����p	��E�����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�(��������V9��V�����%�a��;�6���������l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ہ�����p	��E�����4�
�9�|�w�5��ԜY���F�N��A���;�4��;�%�1��������W9��h��U��%�a��;�6���������l��A�����u�u�u�9�2�W�W���Y���F��1������;�'�9�2�m��������l��R������;�4��9�/����I����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�i�:�������G��h��*���&�2�4�&�0�}����
���l�N��A���;�4��;�%�1��������T9��D��*���6�o�%�:�2�.����4����_%��C��*���y�%�a��9�<�4�������lV��E��U���
�4� �9�8�)����&ù��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�6�(��������V9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��Y��6���'�9�0�e�>�����DӖ��l+��B�����:�
�
�n�w�}�W�������9F�N��U���u�
�
�4�"�1��������9��h��U��%�a��;�6���������l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��<��������_9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�a��;�4��3�����ד�C9��S1��*���
�&�<�;�'�2�W�������@N��1������;�'�9�2�l��������lR��V �����!�:�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�a��;�4��3�����ד�C9��SG�����u�u�u�u�w�}�WϮ�M����F��X �����
�
�%�#�3�4�(���Y����lR��V �����!�:�
�
��-����s���F�R��U���u�u�u�u�w�-�C�������\��X��*ۊ�%�#�1�<��4�W��	�ғ�R��[-�����
�
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ފ�4� �9�:�#�2�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�M����F��X �����
�
�;�&�0�<����&����\��E�����
�
�4� �;�2����&������h#�� ���:�!�:�
������Y����~��V�����9�0�d�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1������;�'�9�2�l�������G��d��U���u�u�u�%�c�����:����\
��h_�����2�i�u�
��<��������_9��UךU���u�u�9�0�]�}�W���Y���C9��z�����;�'�9�0�f�4�(���Y����lR��V �����!�:�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��8���4��;�'�;�8�E���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l+��B�����:�
�
�
�'�+����&����R��P �����o�%�:�0�$�-�C�������\��X��*؊�%�#�1�u����������A	��R1�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l+��B�����:�
�
�
�'�+��������9F�N��U���u�
�
�4�"�1��������9��h��*���&�2�i�u����������A	��R1�����9�n�u�u�w�}����Y���F�N��U���
�4� �9�8�)����&����l��h�����i�u�
�
�6�(��������V9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ǹ��]��t�����0�g�<�
�>�}����Ӗ��P��N����u�
�
�4�"�1��������9��h��*���<�;�%�:�w�}����
�μ�9��Y��6���'�9�0�g�w��(�������]��[1��G���0�y�%�a��3��������l��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�C�������\��X��*؊�%�#�1�|�#�8�W���Y���F���*��� �9�:�!�8��(݁�����Z�G1��8���4��;�'�;�8�E�ԜY���F��D��U���u�u�u�u�'�i�:�������G��h��*���&�2�i�u����������A	��R1�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����4����_%��C��*���
�%�#�1�>�����
������T��[���_�u�u�
��<��������_9��1��*���
�;�&�2�6�.���������T��]���
�4� �9�8�)����&����l��N��A���;�4��;�%�1��������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��<��������_9��1��*���|�u�=�;�]�}�W���Y���C9��z�����;�'�9�0�d�<�(���&����Z�
N��A���;�4��;�%�1��������W]ǻN��U���9�0�_�u�w�}�W���Y����~��V�����9�0�f�4��1�(���
���F��1������;�'�9�2�n��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�a��9�<�4�������lU��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��z�����;�'�9�0�d�4�(���&����T��E��Oʥ�:�0�&�%�c�����:����\
��h]�����;�4��9�/����J����TJ��hZ�����9�:�!�:���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�4� �9�8�)����&����l��G�����_�u�u�u�w�}�W���&����R
��Y�����f�<�
�<�w�`����4����_%��C��*���n�u�u�u�w�8����Y���F�N��*ފ�4� �9�:�#�2�(���&����Z�
N��A���;�4��;�%�1����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�4� �;�2����&����R��[
�����2�4�&�2�w�/����W���F�G1��8���4��;�'�;�8�C���&����Z��^	�����;�%�:�u�w�/����Q����~��V�����9�0�a�4��1�[Ϯ�M����F��X �����
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��8���4��;�'�;�8�C���&����F��R ��U���u�u�u�u�'�i�:�������G��h��*���#�1�<�
�>�}�JϮ�M����F��X �����
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�a��3��������l��h�����<�
�<�u�j�-�C�������\��X��*ފ�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h#�� ���:�!�:�
������Ӈ��Z��G�����u�x�u�u�'�i�:�������G��h��*���&�2�4�&�0�����CӖ��P����*��� �9�:�!�8��(��	�ғ�R��[-�����
�
�
�'�0�}�(ہ�����p	��E�����4�
�9�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����~��V�����9�0�a�4��1�^������F�N��U���%�a��;�6���������l��D��I���
�
�4� �;�2����&����9F�N��U���0�_�u�u�w�}�W���&ǹ��]��t�����0�a�<�
�>�}�JϮ�M����F��X �����
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Y��6���'�9�0�`�6�����������^	�����0�&�u�x�w�}����4����_%��C��*���
�%�#�1�>�����
����l��TN����0�&�%�a��3��������l��h�����u�
�
�4�"�1��������9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����4����_%��C��*���
�%�#�1�~�)����Y���F�N��*ފ�4� �9�:�#�2�(���&����_��Y1����u�
�
�4�"�1��������9��h��N���u�u�u�0�$�}�W���Y���F��hZ�����9�:�!�:���(�������]9��PN�U���
�4� �9�8�)����&ƹ��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������]��[1��@���
�<�u�&�>�3�������KǻN��*ފ�4� �9�:�#�2�(���&����Z��D�����:�u�u�'�4�.�_���&����R
��Y�����`�u�
�
�6�(��������V9��G��Yʥ�a��;�4��3�����ӓ�C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�a��3��������l��h�����|�!�0�u�w�}�W���Y����lR��V �����!�:�
�
��3����E�Ƽ�9��Y��6���'�9�0�`�]�}�W���Y����l�N��U���u�%�a��9�<�4�������lS��Y1����u�
�
�4�"�1��������9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�c�����:����\
��hX�����1�<�
�<�w�.����	����@�CךU���
�
�4� �;�2����&����R��[
�����2�4�&�2��/���	����@��hZ�����9�:�!�:���(������C9��z�����;�'�9�0�a�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�4� �;�2����&����R��[
��U���;�_�u�u�w�}�W���&ǹ��]��t�����0�c�4�
�;��������C9��z�����;�'�9�0�a�<�(���B���F����ߊu�u�u�u�w�}�(ہ�����p	��E�����4�
�9�
�9�.���Y����~��V�����9�0�c�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C�����;�4��9�/����O����@��V�����'�6�&�{�z�W�W���&ǹ��]��t�����0�c�<�
�>���������PF��G�����%�a��;�6���������F��1������;�'�9�2�k����UӖ��l+��B�����:�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hZ�����9�:�!�:���(��������YNךU���u�u�u�u����������A	��R1�����<�u�h�%�c�����:����\
��hX�U���u�u�0�&�w�}�W���Y�����h#�� ���:�!�:�
���������C9��z�����;�'�9�0�a�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*��� �9�:�!�8��(؁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��Y��6���'�9�0�b�6���������l��^	�����u�u�'�6�$�u�(ہ�����p	��E�����4�
�9�y�'�i�:�������G��h��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��Y��6���'�9�0�b�6�����Y����l�N��U���u�%�a��9�<�4�������lQ��G1�����
�<�u�h�'�i�:�������G��h��*���#�1�_�u�w�}�W������F�N��Uʥ�a��;�4��3�����ѓ�C9��S1��*���u�h�%�a��3��������l��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ғ�R��[-�����
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�a��9�<�4�������lQ��Y1�����&�2�
�'�4�g��������lR��V �����!�:�
�
�{�-�C�������\��X��*݊�'�2�u�
��<��������_9�� 1��*���|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ہ�����p	��E�����4�
�9�|�w�5��ԜY���F�N��A���;�4��;�%�1��������TF���*��� �9�:�!�8��(��Y���F��[�����u�u�u�u�w��(�������]��[1��B���
�<�u�h�'�i�:�������G��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�m��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����I����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�G�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*ڊ�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��E�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�e�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�l��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����H����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�F�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*ۊ�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��D�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�d�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�o��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����K����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�E�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*؊�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��G�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�g�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�n��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����J����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�D�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*ي�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��F�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�f�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�i��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����M����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�C�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*ފ�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��A�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�a�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�h��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����L����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�B�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*ߊ�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��@�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�`�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�k��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����O����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�A�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*܊�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��C�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�c�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9�� 1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�j��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����N����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9�� 1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�@�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*݊�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��B�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�b�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�e��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����A����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�O�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*Ҋ�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��M�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�m�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`��;�0�2�d��������l��h�����%�:�u�u�%�>����&ƹ��]��R1�����9�y�%�`��3����@����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����R��[
��U���;�_�u�u�w�}�W���&ƹ��]��R1�����9�
�;�&�0�a�W���&����V9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�4�2�
�
��-��������TF���*���2�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4�2�
������Ӈ��Z��G�����u�x�u�u�'�h�%�������l��D�����2�
�'�6�m�-����
ۖ��l4��P��*���%�`��;�2�8�N�������lS��V ��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��P��*ӊ�%�#�1�|�#�8�W���Y���F���*���2�
�
�
�9�.���Y����a��R1��L�ߊu�u�u�u�;�8�}���Y���F�G1��'���0�0�l�<��4�W��	�ӓ�R��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����^��E��*ڊ�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
�6�<����
����l��A�����<�
�&�<�9�-����Y����V��G1��%���8�!�'�
�������Ƽ�9��E�����
�
�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��C���'�8�!�'���(��������YNךU���u�u�u�u����������l��h�����<�
�<�u�j�-�A�������V��R1�����9�n�u�u�w�}����Y���F�N��U���
�4�4�0�2�.��������W9��h��U��%�c��'�:�)����&ù��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������A��h^�����2�4�&�2�w�/����W���F�G1��%���8�!�'�
����������Z��G��U���'�6�&�}����������l��N��C���'�8�!�'���(����Ƽ�9��E�����
�
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h>�����0�&�0�e�6�����Y����l�N��U���u�%�c��%�0����&����Z��^	��Hʥ�c��'�8�#�/�(���B���F����ߊu�u�u�u�w�}�(ف�����G��h��*���&�2�i�u����������l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������A��h_�����1�<�
�<�w�.����	����@�CךU���
�
�4�4�2�8����H����E
��^ �����&�<�;�%�8�}�W�������C9��g�����'�
�
�
�'�+����&Ź��A��C��*���
�%�#�1�'�8�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����!�'�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�<����
����l��A�����<�u�h�%�a���������V9��V����u�u�u�u�2�.�W���Y���F���*���4�0�0�&�2�l��������l��R������'�8�!�%��(ށ�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��<��������lW��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��g�����'�
�
�
�9�.����
����C��T�����&�}�
�
�6�<����
����F��1�����!�'�
�
��/����&Ź��A��C��*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l6��V�����0�d�4�
�;�t�W������F�N��Uʥ�c��'�8�#�/�(���&����Z�
N��C���'�8�!�'���L���Y�����RNךU���u�u�u�u����������l��h�����i�u�
�
�6�<����
����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��<��������lU��G1�����
�<�u�&�>�3�������KǻN��*܊�4�4�0�0�$�8�D���&����Z��^	�����;�%�:�u�w�/����Q����c��Z�����
�
�%�#�3�}�(ف�����G��h��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��E�����
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�4�4�2�8����J����E
��^ �����h�%�c��%�0����&����R��[
�U���u�u�0�&�w�}�W���Y�����h>�����0�&�0�f�6���������Z�G1��%���8�!�'�
����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�6�8�����Փ�]9��PN�����u�'�6�&�y�p�}���Y����c��Z�����
�
�;�&�0�<����&����\��E�����
�
�4�4�2�8����J�Ƽ�9��E�����
�
�
�'�0�}�(ف�����G��h��*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�O����R��R�����4�
�9�|�w�5��ԜY���F�N��C���'�8�!�'���(���
���F��1�����!�'�
�
�l�}�W���YӃ��VFǻN��U���u�u�
�
�6�<����
����l��D��I���
�
�4�4�2�8����J����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(߁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�e�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(߁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��h^�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ڊ�;�&�2�4�$�:�W�������K��N������<�&�0�g�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����e�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������֓�C9��SG�����u�u�u�u�w�}�WϮ�N����]��h^�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����I����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(ށ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�d�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(ށ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��h_�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ۊ�;�&�2�4�$�:�W�������K��N������<�&�0�f�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����d�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������ד�C9��SG�����u�u�u�u�w�}�WϮ�N����]��h_�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����H����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(݁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�g�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(݁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��h\�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*؊�;�&�2�4�$�:�W�������K��N������<�&�0�e�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����g�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������ԓ�C9��SG�����u�u�u�u�w�}�WϮ�N����]��h\�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����K����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(܁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�f�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(܁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��h]�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ي�;�&�2�4�$�:�W�������K��N������<�&�0�d�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����f�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������Փ�C9��SG�����u�u�u�u�w�}�WϮ�N����]��h]�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����J����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(ہ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�a�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(ہ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��hZ�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ފ�;�&�2�4�$�:�W�������K��N������<�&�0�c�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����a�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������ғ�C9��SG�����u�u�u�u�w�}�WϮ�N����]��hZ�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����M����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(ځ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�`�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(ځ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��h[�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ߊ�;�&�2�4�$�:�W�������K��N������<�&�0�b�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����`�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������ӓ�C9��SG�����u�u�u�u�w�}�WϮ�N����]��h[�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����L����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(ف�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�c�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(ف�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��hX�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*܊�;�&�2�4�$�:�W�������K��N������<�&�0�a�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����c�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������Г�C9��SG�����u�u�u�u�w�}�WϮ�N����]��hX�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����O����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(؁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�b�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(؁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��hY�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*݊�;�&�2�4�$�:�W�������K��N������<�&�0�`�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����b�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������ѓ�C9��SG�����u�u�u�u�w�}�WϮ�N����]��hY�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9�� 1��*���u�h�%�b��4����N����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(ׁ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�m�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(ׁ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��hV�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*Ҋ�;�&�2�4�$�:�W�������K��N������<�&�0�o�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����m�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������ޓ�C9��SG�����u�u�u�u�w�}�WϮ�N����]��hV�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����A����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4�9��(ց�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^ �����4�
�9�
�9�.����
����C��T�����&�}�
�
�6�3�(���&����_�G1��2���&�0�l�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�4�;�
�
��-����PӒ��]FǻN��U���u�u�
�
�6�3�(���&����_��Y1����u�
�
�4�9��(ց�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�R��h��*���#�1�<�
�>�}�JϮ�N����]��hW�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l!��Y��*ӊ�;�&�2�4�$�:�W�������K��N������<�&�0�n�4�(���&����T��E��Oʥ�:�0�&�%�`��������C9��p�����l�%�0�y�'�j�0���
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`������ߓ�C9��SG�����u�u�u�u�w�}�WϮ�N����]��hW�����2�i�u�
��<����&��ƹF�N�����_�u�u�u�w�}�W���&����@9��1��*���u�h�%�b��4����@����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�<�9�1�(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��d�����0�e�4�
�;���������Z��G��U���'�6�&�}����������9��h��Yʥ�l��2�4�$�8�G���&����C��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�>�3����&ù��l��G�����_�u�u�u�w�}�W���&����R
��R1�����9�
�;�&�0�a�W���&����R
��R1�����9�n�u�u�w�}����Y���F�N��U���
�<�;�9���(�������]9��PN�U���
�<�;�9���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�>�3����&ù��l�������%�:�0�&�w�p�W���	�ߓ�Z��[��*ڊ�;�&�2�4�$�:�(�������A	��D��*ӊ�<�;�9�
��q����*����_��h^�����u�
�
�<�9�1�(���&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�<�9�1�(���&����_����ߊu�u�u�u�w�}�(ց�����@9��1��*���u�h�%�l��:��������F�N�����u�u�u�u�w�}�WϮ�@����]��h��*���&�2�i�u����������9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�n�����
����l��A�����<�u�&�<�9�-����
���9F���*���;�9�
�
��-��������T9��D��*���6�o�%�:�2�.����*����_��h_�����1�u�
�
�>�3����&¹��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�d�$�������lW��G1�����!�0�u�u�w�}�W���YӖ��l5��Y��*���
�%�#�1�>�����DӖ��l5��Y��*���
�%�#�1�]�}�W���Y����l�N��U���u�%�l��0�<����H����E
��^ �����h�%�l��0�<����H����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�d�$�������lW��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��d�����0�d�<�
�>���������PF��G�����%�l��2�6�.���Y����`��V�����%�0�y�%�n�����
����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�n�����
����l��A��\ʡ�0�u�u�u�w�}�W���	�ߓ�Z��[��*ۊ�;�&�2�i�w��(�������V9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�
9��P �����d�<�
�<�w�`����*����_��h_�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(ց�����@9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�l��2�4�$�8�E���&����Z��^	�����;�%�:�u�w�/����Q����`��V�����4�
�9�y�'�d�$�������lT��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R
��R1�����9�|�u�=�9�W�W���Y���F��1�����&�0�g�4��1�(���
���F��1�����&�0�g�4��1�L���Y�����RNךU���u�u�u�u����������9��h��*���&�2�i�u����������9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R
��R1�����<�u�&�<�9�-����
���9F���*���;�9�
�
��3��������]9��X��U���6�&�}�
��4����&������h=�����
�
�
�'�0�}�(ց�����@9��1��*���|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ց�����@9��1��*���|�u�=�;�]�}�W���Y���C9��d�����0�g�<�
�>�}�JϮ�@����]��h��N���u�u�u�0�$�}�W���Y���F��hW�����9�
�
�
�9�.���Y����`��V�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����*����_��h\�����'�4�
� �e�o����D������h=�����
�
�
�;�$�:�W������K�d��Uʥ��&�9�
�`�;�(��&���F��G1�����9�d�
�u�w�2�(�������l��d��Uʥ��&�9�
�o�;�(��&���F��h8��G���3�
�g�
�f�n�W������O���*���<�3�
�c��n�L���YӖ��V��C1�*���d�l�
�f�k�}��������_��h^��U���
�
�e�3��m�B���P���F��e�����e�3�
�d�n�-�W��Q����_T��1��*��d�%�}�d�3�*����H���G�� Z��D���
�d�d�%�~�W�W���&����_��1��*��m�%�u�h������A¹��lW��1��]��1�"�!�u�f�}�W���&�ѓ�l ��Z�*��n�u�u�%��.����&���� Q��G]��H���%�6�;�!�;�l�(���Y����e9��h��D��
�a�n�u�w�-�!���&�ߓ�F9��_��D��u�
�d��'�)�(���&����Z��N�����9�
�d�3��o�F���Y����`9��b,�� ���
�0�
�m�a�W�W���&����l��B1�D���u�h�%�d��3�����֓�]9��PUךU���0�
�
�
��i�(�������G9��h_�A���u�h�_�u�w�}�W�������l
��1�Eʢ�0�u�!�%�>�4�ށ�@����U��h�E���u�d�|�0�$�}�W���Y����C9��Y����
�e�n�u�w�/��������
9��D�����3�
�e�`�'�}�J�ԜY���F��h�����#�`�`�e� �8�WǪ�	����l��Q��E���%�}�|�h�p�z�W������F�N��*���&�
�#�`�f�m�}���Y����9��^1�����
�4�!�3��k�(��E��ƹF�N�����;�!�9�d��m�W����θ�C9��^1��FҊ� �m�`�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�B��I���F��C1�����
� �d�g��n�K���Y���F��G1�����9�d�
�e�g�*��������l��1�*���d�d�
�g�g�}�W��PӃ��VFǻN��U���%�6�;�!�;�l�(��I���F��C1�����
� �d�a��n�K���Y���F��G1�����9�d�
�e�g�*��������l��1��*��`�%�}�|�j�z�P������F�N�����:�&�
�#�b�i�G��Y����V��h��*���m�d�%�u�j�W�W���Y�ƭ�l��D�����a�e�u�=�9�u����&���� ^��B1�@���}�|�h�r�p�}����s���F�V�����
�#�`�a�g�f�W���
����^��^Z�� ��b�
�g�i�w�)��������U��\�����:�u�%�6�9�)����H��ƹF��R�����<�
� �d�b��E��Yے��l��h�����f�m�%�u�8�}��������EW��UךU���0�
�8�d�>�;�(��&���F��Z��*���
� �m�l�'�}����	����@��A_��\�ߊu�u�0�
�:�o�ہ�����9��R��]���
�f�
�
��e����I�ߓ�F��SN�����%�
�a�3��m�F���P���F��[1��؊�`�3�
�f�a�-�W��Q����U��^1��ۊ� �d�g�
�e�<�ϭ�����9��h��D���
�g�n�u�w�.����	����U��Y��G��u�!�%�d�f�4��������
9����U���
�8�d�<�1��Oށ�K��ƹF��R�����<�
� �d�`��E��Y���D��F��*����g��!�e�����-����9��h_�F���u�u�%�6�9�)���&����F��D��E��u�u�&�9�#�-�(�������R��N�U��u�=�;�}��%�"�������9��h�����3�
�f�g�'�}�W�������l
��1�E���0�&�u�e�l�}�Wϭ�����9��Q��Mߊ�g�i�u�d�w�5����*����2��x��Gڊ�;�3��%��(�O���	���R��X ��*���`�a�e�|�2�.�W��B�����h��B���
� �d�m��o�K���H�ƻ�V�Q=��8���g��!�g��3����	����U��V�����u�%�6�;�#�1�Fځ�I����_��^�����u�0�
�8�`�4�(���H����CT�
N��Wʢ�0�u�3�
���E����ѓ�]9��c��*���d�c�
�f�j�<�(���
����S��^�����u�e�n�u�w�.����	Ĺ��U��_��G��u�d�u�=�9�u�$���,����|��^������%�
� �o�n����Y����\��h��@��e�u�9�0�u��}���Y����G��h�����d�b�%�u�j�u�����Г�9��h_�@���u�'�&�9�#�-�(�������W��G�U���&�9�!�%��o����M�Г�F�F�����%�
�f�3��i�C���Y����V
��Z��؊� �d�c�
�e�f�W���
����^��^1��*��
�g�i�u�$�1����&����l_��h����0�
�8�b�>�;�(��&���9F���*���
�a�3�
�g�n����D���F�N�����<�<�
� �f�i�(��������h��*���3�
�e�l�'�u�^��^���V
��d��U���u�4�
�:�$�����M����F�D�����<�
� �d�c��D��Y���F���*���
�d�3�
�d�m�������G��^1��ۊ� �d�e�
�e�m�W���H����_��=N��U���u�%�6�;�#�1�Fځ�I��ƹF��R�����
� �m�f�'�}�J�ԜY���F��C1�����3�
�`�
�d�*��������l��h��M���%�}�|�h�p�z�W������F�N��*���&�
�#�`�c�m�}���Y����V��^_�� ��d�
�g�i�w�l�W����ο�T��������;� �
�g�4�(���&����U��W�����i�&�2�0��-��������9��N�����e�n�u�u�#�-�F�������
T��G\��H���w�"�0�u�$�:����*����2��x��Gڊ�;�0�%��f�;�(��&���F��P ��]���6�;�!�9�f��^������D��N�����d�c�3�
�c��F��Y����~3�� ����
�;�0�%��l����Iʹ��^�_�����:�e�n�u�w�)���A����W��h�I����-� ��9�(�(�������C9��1��*��l�%�}�u�w�}�������9F���*��
� �d�d��l�K���*����2��x��B���
�-�
�
��(�F��&���K�
�����e�n�u�u�#�-�F�������U��h�I���d�u�=�;��4��������f*��Y!��*݊�;�0�%��f�;�(��A����Z��^	��´�
�:�&�
�!�e�F�������V�=N��U���
�f�
�
��l����J�ޓ�F�L�U���;�}�:�
��o����K�ғ�F�V�����
�#�
��w�1����[���F��G1�D���<�<�
� �f�i�(��E���F��R ������g�
� �f�l�(��DӇ��P	��C1��M���|�0�&�u�g�f�W������� W��h��*���m�l�%�u�j��Uϩ�����\��h��M���%�u�u�%�4�3����A������RN��W�ߊu�u�8�
�d�;�(��&���FǻN��U���%�6�;�!�;�e�1������G��^1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�m�g�W�W�������l ��_�*��i�u�u�u�w�}��������_��q(�����}�8�
�g�1��F���	����[�I�����u�u�u�u�w�<�(���
����9��=N��U���
�`�3�
�c�m����D���F�N��*���&�
�#�
��*�������� 9��h_�A���}�|�h�r�p�}����s���F�V�����
�#�
�n�w�}����Nǹ��l ��_�*��i�u�!�%�o����M����@��h^�E���<�
� �d�e��D��Y����^��1�����c�
�f�i�w�)���&����U��N����e�
�
�
�"�d�D���P���F��G1�*���l�f�%�u�j�W�W���Y�Ƹ�C9��h��L���%�u�=�;��0�(���@�ѓ�N��S��D���0�&�u�u�w�}�WϪ�	����l ��Z����u�u�!�%�o����HĹ��Z���*���3�
�d�`�'�}�Ϫ�	����l��Q��D���%�|�_�u�w�0�(�������U��N�U���u�u�u�!�'�k�(���H����CU��_��]���
�g�3�
�f�j����P���A�R��U���u�u�u�!�'�l�O���&����l��=N��U���
�a�3�
�d�k����D�θ�C9��h��D��
�g�:�u�:��F؁�&���� _��G\����u�8�
�`�1��C���	���l�N��Uʡ�%�c�
� �f�l�(��������hV�����f�c�%�}�~�`�P���Y����l�N��Uʡ�%�d�e�3��i�O���B�����hV�����
�a�e�%�w�`�_���&�ӓ�F9��\��F��%�e�e�
��o����M�ԓ� O��N�����3�
�g�
�e�a�WǪ�	����F9��1��U���!�%�d�e�>�;�(��&���9F���*���3�
�d�`�'�}�J���[ӑ��]F��^	��³�
���g��)�E߁�����l0��h��D��
�g�u�u�>�3�ǿ�&����G9��V��0���0�&�u�e�l�}�WϪ�	����U��V�����h�w�w�"�2�}�����Ϊ�l��{:��:���b�<�
�-���(���H����CT�	N�����}�%�6�;�#�1�Fׁ�<����_��^�����u�8�
�
�"�d�B���Y���D��_��]���;�1�3�
���E�������Z��O��*ۊ� �l�l�%�~�c�����έ�l��D������|�u�9�2��U�ԜY�Ƹ�C9��^1��*���3�
�f�a�'�}�J���[ӑ��]F��X��*���3�
�f�a�'�}�W�������l
��1�U���0�w�w�_�w�}����&����l ��]�*��i�u�d�u�?�3�_���&����l ��\�*��h�4�
�:�$��ׁ�PӃ��VF�UךU���8�
�
�
�b�;�(��@����[�L�����}�:�
�
�g�;�(��L����F��h�����#�
�|�0�$�}�G��Y����^��h��C���
�e�`�%�w�`�U�������
��h8��D���
�e�`�%�w�}��������ET��G�����w�w�_�u�w�0�(���&����l ��Z�����h�w�w�"�2�}����/����U��[��D��4�
�:�&��+�D��Y����D��d��Uʡ�%�<�<�<�1��Dց�K���W�@��U¹�6��3�
�e��C������]��[��E���9�0�w�w�]�3�W������