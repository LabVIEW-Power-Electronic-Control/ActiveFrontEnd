-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�u� �2�4��������T��_�[���n�_�&�u�2�8��������l��^	��Ĵ�9�_�0�!�#�}�Gݚ�O�Ҋ�lV��h_�����
�
�:�u�$�W�W�������PNǻN��U���u�u�1�<�#�}�W���Y����T��S��C���u�u�u�u�w�}�W������F������u�h�d�n�]�}�W���Y�����h�����u�u�;�0�2�}�J��K���F�d��Uʥ�'�u�_�u�w�}�W�������F�T��ʦ�1�9�2�6�!�>��������W��X����n�_�u�u�w�}�W���Y���F��^ �����:�<�n�_�w�}�W���Y���F�N��U���u�!�
�:�>�����ۂ��W��N�����u�|�_�u�w�}�W�������F�T��ʦ�1�9�2�6�!�>��������W��X����n�_�u�u�w�}�W���Y���F��^ �����:�<�n�_�w�}�W���Y���F�N��U���u�!�
�:�>�����ۂ��W��N�����u�|�_�u�w�}�W������F�N��U���
�:�<�_�w�}�L����Ʃ�G��Nװ���=�!�6� �2�/�ϱ�Y����P��q��*���d�>�'�
��2�W���s����]��V
��E���%�o�&�1�;�:��������R��C��U���;�:�e�n�]�4��������l��T�����:�<�
�0�#�/��������W	��C��\���!�%�u�0��/����
Ӈ��R�N��U���
�<�0�d�w�;��������l��C��]���1�=�d�1� �)�W���Y����]��Z��Oʸ�8�4�'�,�m�}�}���Y�Ƹ�W�L�D��d�d�d�d�f��W���G����W��_�D��d�w�u�u�i��F��H����W��^��U���u�a�h�u�g�l�F��H����W��N�H���e�d�d�d�f�l�G��[����X�_�D��d�d�d�d�u�}�W���N���V��_�D��e�e�e�y�o�`�W��H����W��_�D���l�h�u�e�f�l�F��I����D�=N��U��h�u�e�d�f�l�F��I����F��S�W��d�d�d�e�f�l�F��H���D��_�D��d�e�d�w�w�}�W��Y���W��_�D��d�e�w�u�c�`�W��H����W��^�D���d�u�k�w�f�l�F��H����W�d��U��u�k�w�d�f�l�F��I����J� N��U��d�d�d�e�g�l�F���Y���F�_�D��e�d�e�e�{�W�W���@���V��_�D��e�e�e�y�e�}�I���H����W��^�D���u�d�h�u�g�l�F��H����V��NךU���g�h�u�e�f�l�F��I����D�]��K���d�d�d�e�g�l�G��U����X�_�D��d�e�d�e�u�}�W���K���D��_�D��d�d�d�w�w�k�J���I����W��_�E��y�g�u�k�u�l�F��I����W��B��U���g�u�k�w�f�l�F��I����V�\�H���e�d�d�e�f�l�F��[����[�^�D��d�d�d�d�g�q�}���Y���F�_�D��e�d�e�d�{�n�W���[����W��^�D��w�u�f�h�w�m�F��I����V��L����u�a�h�u�g�l�F��I����W��N�U��w�d�d�d�f�m�G��H���F�L�D��e�d�d�e�g��W���Y����X�_�D��d�d�e�d�u�}�O��Y����W��_�E��d�y�f�u�i��F��H����W��^��U���u�a�u�k�u�l�F��I����V��B��D��u�e�d�d�f�l�F��I���T�	N��D��e�d�d�e�f�m�[�ԜY����[�^�D��d�e�d�e�g�q�C���G����W��_�E��e�w�u�`�j�}�G��H����W��_�Y�ߊu�u�c�h�w�m�F��H����W��L�A���k�w�d�d�g�m�G��H���R��
P��E��d�d�e�d�f�m�U���Y���
F�L�D��d�e�e�e�f��W��D���W��_�E��d�e�y�`�w�c�U��H����W��^�W���u�u�`�u�i��F��I����V��^��U��h�u�e�d�f�m�G��H����F��S�W��d�e�d�e�g�m�G��s���S�	N��D��e�e�d�e�g�m�[��Y���W��^�D��e�e�w�u�`�`�W��H����V��^�E���_�u�u�m�j�}�G��I����W��_�Y���u�k�w�d�f�l�F��H����J�N��U��d�e�d�e�f�l�G���Y���P��
P��E��e�d�e�d�g�l�U���K���V��^�E��d�e�d�y�a�}�I���H����V��^�D���u�u�u�c�w�c�U��H����W��^�W���`�h�u�e�f�m�G��H����D�X��K���d�d�d�d�g�m�F��U���F��S�W��d�d�d�d�f�l�G��O���D��_�E��e�e�e�w�w�d�J���I����V��_�E��y�_�u�u�g�`�W��H����V��^�E���b�u�k�w�f�l�F��I����W�Y�H���e�d�e�d�f�l�G��[��ƹF�N��U��d�e�d�e�g�l�F���Y���F�_�E��e�e�e�e�{�j�W���[����V��^�D��w�u�u�u�`�}�I���H����V��_�E���u�b�h�u�g�l�G��H����W��N�U��w�d�d�e�f�m�F��I���F� W��K���d�d�e�d�f�m�G��U����X�_�E��d�d�e�d�u�}�F��Y����V��_�E��d�y�_�u�w�o�J���I����V��_�E��y�m�u�k�u�l�G��H����V��B��A��u�e�d�d�f�m�G��H���9F�V�H���e�d�d�d�f�l�F��[����[�^�E��e�e�d�d�f�q�O���G����V��^�D��e�w�u�u�w�e�W���[����W��_�D��w�u�l�h�w�m�F��I����V��L�L���k�w�d�e�f�m�F��I���l�N�U��w�d�e�d�g�m�G��H���F�L�D��e�e�d�e�g��W��D���W��_�E��e�e�y�_�w�}�C��Y����W��^�E��d�y�l�u�i��F��I����W��_��U��h�u�e�d�f�l�G��H����FǻN��B��u�e�d�d�g�l�F��I���
^�	N��D��e�d�e�e�f�m�[��Y���W��^�E��d�d�w�u�w�}�F��D���W��^�E��d�d�y�d�f�`�W��H����V��^�E���d�g�h�u�g�l�G��H����V��NךU���e�u�k�w�f�m�F��H����W�_�U��w�d�e�d�g�l�F��I���S�	N��D��d�e�d�d�f�l�[�ԜY����F�L�D��e�d�e�d�f��W��Y���W��_�E��e�e�w�u�g�}�I���H����V��^�E���u�u�u�d�n�`�W��H����V��_�E���d�e�h�u�g�l�G��H����W��N�D��u�e�d�e�f�m�F��I���9F�_�U��w�d�e�e�g�l�F��I���U�	N��D��e�e�d�d�g�m�[��M���V��^�D��d�e�d�y�]�}�W��Y���W��^�E��d�d�w�u�f�}�I���H����V��^�E���u�d�u�k�u�l�G��I����V��B��U���d�m�h�u�g�m�F��H����V��N�L��u�e�e�d�f�m�G��H���T��
P��E��d�d�d�e�g�l�U���Y���W�	N��D��d�e�d�d�g�m�[��K���V��_�D��e�e�e�y�f�n�J���I����V��_�D��y�_�u�u�e�}�I���H����V��_�E���u�g�u�k�u�l�F��I����V��B��G���k�w�d�d�g�l�G��H���l�N�B��u�e�e�d�f�m�G��I���T��
P��E��d�d�d�e�g�l�U���K���D��_�E��d�e�e�w�w�}�W��I���V��_�D��e�d�e�y�f�l�J���I����V��^�D��y�d�g�h�w�m�G��I����V��L����u�f�u�k�u�l�F��H����V��B��F���k�w�d�d�f�l�G��H���W��S�W��d�d�e�e�g�m�G��s���U��
P��E��e�e�d�d�g�l�U���J���D��_�E��d�e�e�w�w�n�W���[����W��_�D��w�u�u�u�f�d�J���I����V��_�E��y�d�e�h�w�m�G��H����W��L�D��h�u�e�e�g�l�G��I����FǻN��A���k�w�d�d�g�m�F��I���W��S�W��d�e�d�d�g�l�F��H���F�^�E��e�d�d�e�{�W�W���M���D��_�E��e�d�e�w�w�i�W���[����W��_�D��w�u�a�u�i��F��H����W��^��U���u�d�m�h�w�m�G��H����V��L�D��h�u�e�e�f�l�G��I����F��N��U��e�d�e�d�g�m�G���Y���W��S�W��e�d�e�d�g�m�F��H���F�^�D��d�e�e�e�{�l�D��Y����W��_�D��e�y�_�u�w�h�W���[����V��_�D��w�u�`�u�i��F��I����W��^��U���u�k�w�d�g�m�F��H����J�N��D��h�u�e�e�f�m�G��H����F��N��U��e�d�e�e�f�l�F���Y����X�_�E��d�e�e�e�u�}�W���H���F�^�D��e�d�d�d�{�l�F��Y����V��^�D��d�y�d�g�j�}�G��I����V��^�Y�ߊu�u�c�u�i��F��H����V��^��U��u�k�w�d�g�l�G��H����J�[��K���d�e�e�d�f�l�G��U���F��N��U��e�e�d�e�f�m�F���Y����X�_�E��e�d�d�d�u�}�A���G����V��_�E��d�w�u�u�w�l�N��Y����V��^�E��d�y�d�e�j�}�G��I����W��^�Y��d�h�u�e�f�l�F��I����D�=N��U��u�k�w�e�f�l�F��H����J� ]��K���e�d�d�e�f�m�G��U����[�^�D��d�e�d�e�g�q�}���Y����X�^�D��e�e�d�e�u�}�@���G����W��^�E��d�w�u�b�w�c�U��H����V��_�W���u�u�d�m�j�}�G��H����W��_�Y��l�h�u�e�f�l�F��I����D�V�H���e�d�d�e�f�m�F��[��ƹF�_��K���e�d�e�e�f�l�G��U����[�^�D��e�e�e�d�f�q�F��D���W��_�D��e�e�y�_�w�}�O���G����W��^�D��d�w�u�m�w�c�U��H����V��_�W���m�u�k�w�g�l�F��H����V�d��U��b�h�u�e�f�m�G��I����D�V�H���e�d�e�d�f�m�F��[����
F�L�D��d�e�d�e�f��W���Y����[�^�D��e�d�e�d�g�q�F��D���W��^�E��d�d�y�d�e�`�W��H����W��_�E���_�u�u�l�w�c�U��H����W��^�W���l�u�k�w�g�m�F��I����W�_�U��w�e�e�d�g�l�G��I���F�W�H���e�d�d�d�g�m�G��[����F�L�D��e�e�e�e�g��W��Y���V��_�D��d�e�w�u�w�}�F��D���W��_�D��d�e�y�g�g�`�W��H����V��_�D���g�d�h�u�g�l�F��I����W��NךU���e�u�k�w�g�m�G��I����V�\�U��w�e�e�e�g�l�G��H���R�	N��E��e�e�e�e�f�l�[�ԜY����F�L�D��d�e�d�d�g��W��Y���V��_�D��d�e�w�u�g�}�I���I����W��^�E���u�u�u�g�o�`�W��H����V��_�E���g�l�h�u�g�l�G��I����W��N�E��u�e�d�e�f�l�F��H���9F�\�U��w�e�e�e�g�l�G��H���T�	N��E��e�e�e�e�f�m�[��J���V��^�D��e�e�e�y�]�}�W��Y���V��^�D��d�d�w�u�f�}�I���I����W��_�E���u�d�u�k�u�m�F��H����V��B��U���g�b�h�u�g�m�F��I����W��N�M��u�e�e�d�g�l�G��H���W��
P��E��d�e�d�e�g�m�U���Y���V�	N��E��d�e�e�e�f�m�[��H���V��_�D��e�d�d�y�e�o�J���I����W��^�E��y�_�u�u�e�}�I���I����W��_�D���u�g�u�k�u�m�F��I����V��B��G���k�w�e�d�g�m�G��I���l�N�C��u�e�e�e�f�m�F��H���T��
P��E��e�d�d�d�f�m�U���K���D��_�E��d�e�d�w�w�}�W��@���V��^�D��d�d�e�y�e�m�J���I����V��^�D��y�g�d�h�w�m�G��H����W��L����u�f�u�k�u�m�F��I����V��B��F���k�w�e�d�g�m�G��I���T��S�W��d�e�d�e�f�m�G��s���U��
P��E��e�e�e�d�g�l�U���J���D��^�D��d�d�d�w�w�n�W���[����W��_�E��w�u�u�u�e�e�J���I����W��^�D��y�g�l�h�w�m�G��I����V��L�G��h�u�e�e�f�m�F��H����FǻN��A���k�w�e�e�g�l�F��H���T��S�W��e�e�e�d�f�m�F��K���F�^�E��e�d�e�d�{�W�W���M���D��^�E��d�d�d�w�w�i�W���[����V��^�E��w�u�a�u�i��G��H����W��_��U���u�g�b�h�w�m�G��H����V��L�G��h�u�e�e�g�l�G��H����F��N��U��e�e�e�e�f�l�F���Y���T��S�W��e�d�e�e�f�l�G��K���F�^�E��d�e�d�d�{�o�E��Y����V��^�E��e�y�_�u�w�h�W���[����V��_�D��w�u�`�u�i��G��I����W��^��U���u�k�w�e�g�m�G��I����J�N��G��h�u�e�e�g�m�G��I����F�� N��U��d�d�d�e�f�m�F���Y����X�_�D��e�d�d�d�u�}�W���K���F�_�D��e�e�d�d�{�o�G��Y����W��_�D��e�y�g�d�j�}�F��H����V��_�Y�ߊu�u�c�u�i��F��I����V��^��U��u�k�w�d�f�m�G��I����J�Z��K���d�d�e�d�g�l�G��U���F��N��U��d�d�e�d�f�l�F���Y����X�_�D��e�d�e�d�u�}�A���G����W��_�E��d�w�u�u�w�o�O��Y����V��_�D��d�y�g�l�j�}�F��I����V��^�Y��e�h�u�d�f�m�G��I����D�=N��U��u�k�w�d�f�l�G��H����J� \��K���d�d�e�d�f�l�F��U����[�_�D��e�e�e�d�g�q�}���Y����X�_�E��d�d�e�e�u�}�@���G����W��_�E��e�w�u�b�w�c�U��H����W��_�W���u�u�g�b�j�}�F��H����V��^�Y��m�h�u�d�f�l�F��I����D�Y�H���d�d�d�e�f�l�F��[��ƹF�^��K���d�e�d�d�g�l�G��U����[�_�E��e�d�d�e�f�q�E��D���W��_�E��e�d�y�_�w�}�O���G����V��^�D��e�w�u�m�w�c�U��I����V��_�W���m�u�k�w�f�m�G��H����V�d��U��c�h�u�d�f�l�G��I����D�V�H���d�d�e�d�f�m�F��[����F�L�D��d�e�e�e�f��W���Y����[�_�E��e�d�e�e�g�q�E��D���W��^�D��d�d�y�g�f�`�W��H����W��_�D���_�u�u�l�w�c�U��I����W��_�W���l�u�k�w�f�m�G��I����V�\�U��w�d�e�e�g�l�G��H���F�W�H���d�d�e�e�f�l�F��[����F�L�D��e�d�d�e�f��W��Y���W��^�E��e�d�w�u�w�}�E��D���V��_�D��e�d�y�g�n�`�W��I����W��_�E���f�e�h�u�f�m�F��H����V��NךU���e�u�k�w�f�l�F��I����W�]�U��w�d�d�d�g�l�F��H���U�	N��D��e�d�e�d�g�l�[�ԜY����F�L�E��d�d�e�d�g��W��Y���W��^�E��d�e�w�u�g�}�I���H����W��_�E���u�u�u�f�`�`�W��I����W��_�E���f�m�h�u�f�m�G��H����V��N�L��u�d�e�e�f�m�G��H���9F�]�U��w�d�d�d�g�l�F��I���W�	N��D��d�d�e�d�f�m�[��K���W��^�E��e�e�d�y�]�}�W��Y���W��_�E��e�e�w�u�f�}�I���H����W��^�D���u�d�u�k�u�l�F��I����V��B��U���f�c�h�u�f�m�G��H����W��N�B��u�d�e�e�g�m�F��I��� W��
P��D��e�e�e�d�f�m�U���Y���_�	N��D��d�d�e�d�f�m�[��I���W��_�D��e�d�e�y�d�l�J���H����W��^�E��y�_�u�u�e�}�I���H����W��_�D���u�g�u�k�u�l�G��I����V��B��G���k�w�d�e�f�m�G��I���l�N�@��u�d�e�d�f�m�F��I��� T��
P��D��d�d�d�d�g�l�U���K���D��^�E��d�d�e�w�w�}�W��A���W��_�D��e�d�e�y�d�d�J���H����V��^�E��y�f�e�h�w�l�G��H����W��L����u�f�u�k�u�l�G��H����W��B��F���k�w�d�e�f�m�F��I���U��S�W��e�d�d�d�g�m�G��s��� U��
P��D��e�e�e�e�f�m�U���J���D��^�E��e�d�d�w�w�n�W���[����V��^�D��w�u�u�u�d�j�J���H����W��_�E��y�f�m�h�w�l�G��H����W��L�F��h�u�d�e�g�m�F��H����FǻN��A���k�w�d�e�g�m�F��I���U��S�W��e�e�e�e�f�m�G��J���F�_�D��e�e�d�e�{�W�W���M���D��_�D��e�d�d�w�w�i�W���[����W��^�E��w�u�a�u�i��G��H����V��^��U���u�f�c�h�w�l�F��I����W��L�F��h�u�d�d�f�m�G��H����F��N��U��d�d�d�d�g�m�G���Y���U��S�W��d�e�e�d�f�l�G��J���F�_�E��e�d�e�d�{�n�F��Y����W��_�E��d�y�_�u�w�h�W���[����V��_�E��w�u�`�u�i��G��I����W��^��U���u�k�w�e�f�l�F��H����J�N��F���h�u�d�d�g�l�F��I����F��N��U��d�e�d�e�g�l�G���Y����X�^�E��d�d�d�e�u�}�W���J���F�_�D��e�e�d�d�{�n�N��Y����V��^�E��e�y�f�e�j�}�F��I����V��^�Y�ߊu�u�c�u�i��G��I����W��_��U��u�k�w�e�f�m�G��H����J�]��K���e�d�e�d�f�l�F��U���F��N��U��d�e�e�e�g�m�G���Y����X�^�E��d�d�e�d�u�}�A���G����W��^�E��e�w�u�u�w�n�@��Y����W��^�E��e�y�f�m�j�}�F��H����V��^�Y��l�h�u�d�f�l�F��H����D�=N��U��u�k�w�e�g�l�F��H����J� _��K���e�e�d�e�f�l�F��U����[�_�E��e�d�e�d�f�q�}���Y����X�^�D��d�e�d�e�u�}�@���G����V��_�D��d�w�u�b�w�c�U��I����V��^�W���u�u�f�c�j�}�F��H����V��_�Y��b�h�u�d�f�l�G��H����D�Y�H���d�d�d�e�f�l�G��[��ƹF� W��K���e�e�e�e�f�m�F��U����[�_�E��d�e�d�d�f�q�D��D���W��_�E��d�e�y�_�w�}�O���G����V��^�E��e�w�u�m�w�c�U��I����V��_�W���m�u�k�w�g�m�F��H����V�d��U��`�h�u�d�f�m�G��H����D�V�H���d�d�e�e�g�l�G��[����F�L�D��d�d�e�e�f��W���Y����[�_�E��d�d�e�d�g�q�D��D���W��_�D��e�e�y�f�g�`�W��H����V��_�E���_�u�u�l�w�c�U��I����V��^�W���l�u�k�w�g�m�G��I����W�]�U��w�e�e�e�g�m�G��I���F�W�H���d�d�e�e�g�m�F��[����F�L�E��d�d�e�d�g��W��Y���V��_�E��e�e�w�u�w�}�D��D���V��_�E��e�d�y�f�o�`�W��I����V��_�D���f�l�h�u�f�m�F��H����W��NךU���e�u�k�w�g�l�F��I����V�Z�U��w�e�d�d�g�m�G��H���T�	N��E��d�e�e�d�g�l�[�ԜY���� F�L�E��d�d�e�e�g��W��Y���V��^�E��e�d�w�u�g�}�I���I����V��_�E���u�u�u�a�a�`�W��I����V��^�E���a�b�h�u�f�m�F��H����V��N�M��u�d�e�d�g�m�F��I���9F�Z�U��w�e�d�e�g�m�F��H���V�	N��E��e�e�d�e�g�l�[��H���W��^�D��e�d�e�y�]�}�W��Y���V��_�E��d�e�w�u�f�}�I���I����V��^�D���u�d�u�k�u�m�F��I����W��B��U���a�`�h�u�f�m�G��I����W��N�C��u�d�e�e�g�l�G��H���W��
P��D��e�e�e�d�g�l�U���Y���^�	N��E��d�e�e�d�f�l�[��@���W��^�E��e�e�e�y�c�m�J���H����W��^�D��y�_�u�u�e�}�I���I����W��_�E���u�g�u�k�u�m�F��H����W��B��G���k�w�e�d�g�m�G��H���l�N�A��u�d�e�e�f�m�F��H���T��
P��D��e�e�d�e�f�l�U���K���D��_�E��d�d�e�w�w�}�W��N���W��^�D��e�d�d�y�c�e�J���H����V��_�E��y�a�l�h�w�l�G��I����W��L����u�f�u�k�u�m�G��H����W��B��F���k�w�e�e�f�l�F��H���R��S�W��e�d�d�e�f�l�F��s���U��
P��D��d�d�d�d�f�l�U���J���D��^�D��d�e�d�w�w�n�W���[����W��^�E��w�u�u�u�c�k�J���H����V��_�E��y�a�b�h�w�l�G��I����V��L�A��h�u�d�e�f�m�F��H����FǻN��F���k�w�e�e�f�m�G��I���R��S�W��e�d�e�d�g�m�G��M���F�^�E��d�d�d�d�{�W�W���M���D��^�D��d�e�e�w�w�i�W���[����V��_�D��w�u�a�u�i��G��I����W��_��U���u�a�`�h�w�l�G��H����W��L�A��h�u�d�e�f�l�G��H����F�� N��U��e�d�d�e�g�l�G���Y���R��S�W��e�e�d�e�f�l�G��M���F�^�E��d�d�e�e�{�i�G��Y����W��^�E��d�y�_�u�w�h�W���[����V��_�D��w�u�`�u�i��G��I����W��^��U���u�k�w�e�g�m�G��I����J�N��A��h�u�d�e�f�m�G��I����F��N��U��e�e�d�d�g�m�G���Y����X�^�E��e�d�d�d�u�}�W���M���F�^�D��e�d�e�e�{�i�O��Y����V��_�D��e�y�a�l�j�}�F��I����W��_�Y�ߊu�u�c�u�i��G��H����W��^��U��u�k�w�e�g�l�G��H����J�\��K���e�e�d�d�f�l�G��U���F��N��U��e�e�e�d�f�l�F���Y����X�^�E��d�e�e�d�u�}�A���G����V��_�E��e�w�u�u�w�i�A��Y����V��^�D��d�y�a�b�j�}�F��I����V��^�Y��m�h�u�d�g�m�G��H����D�=N��U��u�k�w�e�g�l�G��I����J� ^��K���e�e�d�e�g�l�G��U����[�_�E��e�e�e�d�f�q�}���Y����X�^�E��d�e�e�d�u�}�@���G����V��_�D��d�w�u�b�w�c�U��I����W��_�W���u�u�a�`�j�}�F��I����V��^�Y��c�h�u�d�g�m�F��I����D�Y�H���d�e�e�d�f�l�G��[��ƹF� V��K���e�e�e�e�f�m�F��U����[�_�E��e�e�d�d�f�q�C��D���V��_�D��d�e�y�_�w�}�O���G����V��^�E��d�w�u�m�w�c�U��I����V��^�W���m�u�k�w�g�m�G��I����W�d��U��a�h�u�d�g�m�G��H����D�V�H���d�e�e�e�f�m�G��[����F�L�E��e�d�d�e�g��W���Y����[�_�E��d�e�e�e�f�q�C��D���V��^�D��e�d�y�a�n�`�W��I����V��^�E���_�u�u�l�w�c�U��I����V��^�W���l�u�k�w�g�m�G��I����V�Z�U��w�e�e�e�g�l�F��I���F�W�H���d�e�e�e�f�m�F��[����F�L�E��e�d�e�d�g��W��Y���V��^�D��e�d�w�u�w�}�C��D���V��^�E��d�e�y�a�`�`�W��I����W��_�D���a�m�h�u�f�m�G��I����V��NךU���l�u�k�w�g�m�G��H����V�[�U��w�e�e�e�g�l�F��H���W�	N��E��e�e�d�e�g�l�[�ԜY����F�L�E��e�e�d�d�f��W��Y���V��^�E��e�d�w�u�g�}�I���I����V��^�D���u�u�u�`�b�`�W��I����V��_�E���`�c�h�u�f�m�G��I����W��N�B��u�d�e�e�g�m�G��H���9F�[�U��w�e�e�e�g�m�G��I���_�	N��E��e�e�e�e�f�m�[��I���W��^�E��e�e�e�y�]�}�W��Y���V��^�E��e�e�w�u�f�}�I���I����V��^�E���u�d�u�k�u�m�G��I����V��B��U���`�a�h�u�f�m�G��I����W��N�@��u�d�e�e�g�m�G��H���W��
P��D��e�e�e�e�f�l�U���Y���Q�	N��E��e�e�e�e�f�l�[��A���W��^�E��d�d�e�y�b�d�J���H����V��^�D��y�_�u�u�e�}�I���I����V��^�D���u�g�u�k�u�m�G��I����V��B��G���k�w�e�e�g�m�G��H���l�N�F��u�d�e�e�g�m�G��H���T��
P��D��e�e�e�e�f�m�U���K���D��^�E��d�d�e�w�w�}�W��O���W��^�E��d�e�d�y�b�j�J���H����V��^�E��y�`�m�h�w�l�G��I����W��L����u�g�u�k�u�m�G��I����V��B��F���k�w�e�e�g�m�F��I���S��S�W��e�e�e�d�f�l�G��s���U��
P��D��e�e�d�d�g�l�U���J���D��^�E��e�e�e�w�w�n�W���[����V��^�D��w�u�u�u�b�h�J���H����V��^�D��y�`�c�h�w�l�G��I����V��L�@��h�u�d�e�g�m�F��I����FǻN��F���k�w�e�e�g�l�G��I���S��S�W��e�e�d�d�g�m�F��L���F�^�E��d�e�e�e�{�W�W���M���D��^�D��e�e�e�w�w�i�W���[����V��^�D��w�u�a�u�i��G��I����V��_��U���u�`�a�h�w�l�G��H����V��L�@���h�u�d�e�g�l�F��H����F��N��U��e�e�d�d�g�m�F���Y���S��S�W��e�e�e�d�f�m�F��L���F�^�E��e�d�d�e�{�h�N��Y����V��^�E��d�y�_�u�w�h�W���[����V��_�E��w�u�`�u�i��G��I����V��^��U���u�k�w�e�g�m�F��H����J�N��@��h�u�d�e�g�m�G��I����F��N��U��e�e�e�e�f�l�F���Y����X�^�E��e�d�d�d�u�}�W���L���F�^�D��e�e�e�d�{�h�@��Y����V��_�D��d�y�`�m�j�}�F��I����V��^�Y�ߊu�u�`�u�i��G��H����V��_��U��u�k�w�e�g�l�F��I����J�_��K���e�e�d�d�g�l�F��U���F��N��U��e�e�e�d�f�l�F���Y����X�^�E��e�d�e�d�u�}�A���G����V��^�D��d�w�u�u�w�h�B��Y����V��_�D��e�y�`�c�j�}�F��I����W��_�Y���b�h�u�d�g�m�F��H����D�=N��U��u�k�w�e�g�l�F��H����J�W��K���e�e�d�d�f�m�G��U����[�_�E��e�e�e�d�f�q�}���Y����X�^�D��e�e�d�e�u�}�@���G����V��^�E��e�w�u�b�w�c�U��I����W��_�W���u�u�`�a�j�}�F��H����W��_�Y���`�h�u�d�g�l�G��H����D�Y�H���d�e�d�e�f�l�F��[��ƹF� Y��K���e�e�e�e�g�m�F��U����[�_�E��e�d�d�e�g�q�B��D���V��_�E��e�e�y�_�w�}�O���G����V��^�D��d�w�u�m�w�c�U��I����W��_�W���m�u�k�w�g�m�G��I����V�d��U���f�h�u�d�g�l�F��H����D�V�H���d�e�d�e�g�m�F��[����F�L�E��e�d�d�e�g��W���Y����[�_�E��e�d�d�e�g�q�B��D���V��^�D��e�d�y�`�o�`�W��I����W��_�D���_�u�u�m�w�c�U��I����V��_�W���l�u�k�w�g�m�F��H����V�[�U��w�e�e�d�g�m�F��H���F�W�H���d�e�d�d�g�m�F��[���� F�L�E��d�e�d�d�g��W��Y���V��_�D��d�e�w�u�w�}�B��D���V��^�E��d�e�y�`�a�`�W��I����W��^�D���`�b�h�u�f�m�G��I����V��NךU���l�u�k�w�g�l�G��H����W�[�U��w�e�d�e�f�l�G��H���V�	N��E��e�e�e�d�f�m�[�ԜY����F�L�E��d�d�e�d�f��W��Y���V��^�E��e�d�w�u�g�}�I���I����W��_�E���u�u�u�c�c�`�W��I����W��_�E���c�`�h�u�f�m�G��I����V��N�C��u�d�e�e�g�l�F��I���9F�X�U��w�e�d�d�f�m�G��H���^�	N��E��d�d�e�d�g�m�[��@���W��^�E��e�e�d�y�]�}�W��Y���V��_�E��e�e�w�u�f�}�I���I����V��^�D���u�d�u�k�u�m�F��H����V��B��U���c�f�h�u�f�m�G��H����W��N�A��u�d�e�d�g�m�G��H���W��
P��D��d�e�d�d�f�m�U���Y���P�	N��E��e�d�e�d�g�m�[��N���W��_�D��e�e�d�y�a�e�J���H����W��_�E��y�_�u�u�f�}�I���I����V��_�E���u�g�u�k�u�m�F��H����W��B��G���k�w�e�d�g�l�G��H���l�N�G��u�d�e�d�g�m�G��I���T��
P��D��d�e�d�e�f�l�U���K���D��_�E��e�d�d�w�w�}�W��L���W��_�D��e�d�e�y�a�k�J���H����W��^�D��y�c�b�h�w�l�G��H����V��L����u�g�u�k�u�m�F��H����W��B��G���k�w�e�d�f�l�G��I���P��S�W��e�e�e�e�f�l�G��s���U��
P��D��e�e�d�d�g�l�U���J���D��^�E��d�d�e�w�w�n�W���[����V��^�E��w�u�u�u�a�i�J���H����W��_�E��y�c�`�h�w�l�F��H����V��L�C��h�u�d�d�g�l�G��H����FǻN��F���k�w�e�e�g�l�F��H���P��S�W��e�d�e�d�g�m�F��O���F�_�D��d�d�e�e�{�W�W���M���D��^�E��d�d�d�w�w�i�W���[����W��^�D��w�u�a�u�i��G��H����W��^��U���u�c�f�h�w�l�F��H����W��L�C��h�u�d�d�g�l�F��H����F��N��U��d�d�e�e�g�l�F���Y���P��S�W��e�e�e�d�g�m�G��O���F�_�E��d�d�d�e�{�k�O��Y����W��^�E��e�y�_�u�w�i�W���[����V��^�E��w�u�`�u�i��G��I����W��^��U���u�k�w�e�g�m�F��I����J�N��C��h�u�d�d�f�m�G��I����F��N��U��d�d�e�d�f�l�G���Y����X�^�D��d�e�e�d�u�}�W���O���F�_�D��e�d�e�d�{�k�A��Y����W��_�E��e�y�c�b�j�}�F��H����W��^�Y�ߊu�u�`�u�i��G��I����V��_��U���u�k�w�e�f�m�G��I����J�^��K���e�d�e�d�f�m�G��U���F��N��U��d�e�e�d�g�l�F���Y����X�^�E��e�d�d�d�u�}�A���G����W��_�E��d�w�u�u�w�k�C��Y����V��_�E��e�y�c�`�j�}�F��I����W��_�Y��c�h�u�d�f�m�G��I����D�=N��U��u�k�w�e�f�l�F��I����J�V��K���e�d�d�e�f�m�F��U����[�_�D��e�d�d�e�f�q�}���Y����X�^�E��d�e�e�d�u�}�@���G����W��^�D��e�w�u�b�w�c�U��H����W��^�W���u�u�c�f�j�}�F��H����V��_�Y��a�h�u�d�f�l�F��H����D�Y�H���d�d�d�d�f�m�F��[��ƹF� X��K���e�d�e�d�g�m�F��U����[�_�D��e�e�e�d�f�q�A��D���W��^�D��e�e�y�_�w�}�@���G����W��_�E��d�w�u�m�w�c�U��H����V��^�W���m�u�k�w�g�l�F��H����W�d��U��g�h�u�d�f�l�F��I����D�V�H���d�e�e�e�g�l�F��[����F�L�E��e�d�d�d�g��W���Y����[�_�E��d�e�d�e�g�q�A��D���V��_�D��e�e�y�c�`�`�W��I����W��_�E���_�u�u�m�w�c�U��I����V��^�W���m�u�k�w�f�m�F��H����W�X�U��w�d�e�d�f�m�G��H���F�W�H���d�e�e�e�f�m�G��[����F�L�E��d�e�d�e�f��W��Y���W��_�E��e�d�w�u�w�}�A��D���V��_�D��e�d�y�c�b�`�W��I����W��^�E���c�c�h�u�f�m�F��I����W��NךU���l�u�k�w�f�m�G��H����V�X�U��w�d�e�e�g�m�F��I���
_�	N��D��e�d�d�e�g�l�[�ԜY����F�L�E��e�e�d�e�g��W��Y���W��_�D��d�e�w�u�g�}�I���H����W��_�D���u�u�u�b�d�`�W��I����V��_�D���b�a�h�u�f�m�F��I����V��N�@��u�d�e�d�f�l�F��H���9F�Y�U��w�d�d�e�g�l�F��H���Q�	N��D��e�d�e�d�f�m�[��A���W��^�D��e�d�d�y�]�}�W��Y���W��^�D��d�d�w�u�f�}�I���H����W��^�D���u�d�u�k�u�l�F��I����W��B��U���b�g�h�u�f�m�G��H����V��N�F��u�d�e�e�g�l�G��H���W��
P��D��e�d�e�e�f�m�U���Y���S�	N��D��d�d�e�d�g�l�[��O���W��^�D��d�e�d�y�`�j�J���H����V��^�E��y�_�u�u�f�}�I���H����W��_�E���u�d�u�k�u�l�F��I����V��B��G���k�w�d�d�g�m�F��I���l�N�D��u�d�e�d�f�l�G��I���T��
P��D��d�e�e�e�f�m�U���K���D��_�E��e�d�d�w�w�}�W��M���W��_�D��d�d�e�y�`�h�J���H����W��^�D��y�b�c�h�w�l�G��H����V��L����u�g�u�k�u�l�G��I����V��B��G���k�w�d�e�g�m�F��H���Q��S�W��e�e�d�e�g�m�F��s���U��
P��D��e�d�e�d�f�m�U���J���D��^�D��d�e�e�w�w�n�W���[����V��_�E��w�u�u�u�`�n�J���H����V��_�E��y�b�a�h�w�l�F��I����W��L�B���h�u�d�d�g�l�G��I����FǻN��F���k�w�d�e�f�l�G��H���Q��S�W��e�d�d�d�g�l�F��N���F�_�E��e�d�e�e�{�W�W���J���D��^�E��e�d�e�w�w�i�W���[����V��^�D��w�u�a�u�i��F��I����V��^��U���u�b�g�h�w�l�F��H����W��L�B��h�u�d�d�f�m�G��I����F��N��U��d�d�e�e�f�l�G���Y���Q��S�W��e�d�d�d�f�l�F��N���F�_�D��d�e�d�e�{�j�@��Y����W��_�E��d�y�_�u�w�i�W���[����V��_�E��w�u�a�u�i��F��I����W��^��U���u�k�w�d�f�m�F��I����J�N��B��h�u�d�d�g�l�F��H����F��N��U��d�e�d�e�f�m�G���Y����X�_�E��e�d�d�e�u�}�W���N���F�_�D��e�e�d�d�{�j�B��Y����V��_�E��d�y�b�c�j�}�F��I����V��^�Y�ߊu�u�`�u�i��F��H����W��^��U���u�k�w�d�f�m�G��I����J�W��K���d�d�e�e�f�m�F��U���F��N��U��d�d�e�d�f�l�G���Y����X�_�D��d�e�e�e�u�}�A���G����W��_�E��d�w�u�u�w�j�D��Y����W��^�D��d�y�b�a�j�}�F��H����V��^�Y��`�h�u�d�f�l�G��H����D�=N��U��u�k�w�d�f�l�G��I����J�Y��K���d�d�d�d�g�l�F��U����[�^�E��e�e�e�e�g�q�}���Y����X�^�E��d�e�d�e�u�}�@���G����V��_�E��d�w�u�b�w�c�U��I����W��^�W���u�u�b�g�j�}�G��I����W��^�Y��f�h�u�e�g�m�F��H����D� Y�H���e�e�e�e�f�l�G��[��ƹF� [��K���e�e�d�d�f�l�F��U����[�^�E��e�d�e�e�g�q�@��D���V��_�E��e�d�y�_�w�}�@���G����V��_�E��e�w�u�b�w�c�U��I����V��^�W���m�u�k�w�g�m�G��H����W�d��U��d�h�u�e�g�l�F��H����D� V�H���e�e�d�d�f�l�F��[���� F�L�E��d�d�e�e�g��W���Y����[�^�E��e�e�e�d�g�q�@��D���V��^�D��d�e�y�b�a�`�W��I����V��_�E���_�u�u�m�w�c�U��I����W��_�W���m�u�k�w�g�m�F��I����W�Y�U��w�e�d�e�g�l�F��H���F� W�H���e�e�e�e�g�l�F��[����F�L�E��d�e�e�e�g��W��Y���V��^�D��d�e�w�u�w�}�@��D���V��_�E��d�d�y�b�c�`�W��I����V��^�D���b�`�h�u�g�m�G��I����V��NךU���l�u�k�w�g�l�F��H����V�Y�U��w�e�d�d�g�m�G��I���
^�	N��E��d�d�d�e�f�m�[�ԜY����
F�L�E��e�e�d�e�f��W��Y���V��^�D��d�e�w�u�g�}�I���I����W��_�D���u�u�u�m�e�`�W��I����W��^�D���m�f�h�u�g�m�F��I����W��N�A��u�e�e�d�g�m�G��I���9F�V�U��w�e�d�d�g�l�F��I���P�	N��E��d�d�e�d�g�l�[��N���V��_�E��d�d�d�y�]�}�W��Y���V��_�E��d�d�w�u�g�}�I���I����W��_�E���u�d�u�k�u�m�G��I����W��B��U���m�d�h�u�g�l�G��I����W��N�G��u�e�d�e�f�m�F��I���W��
P��E��e�d�d�d�g�m�U���Y���R�	N��E��e�d�e�e�f�l�[��L���V��^�E��e�d�d�y�o�k�J���I����V��_�E��y�_�u�u�f�}�I���I����W��^�E���u�d�u�k�u�m�G��I����V��B��D���k�w�e�e�f�l�F��I���l�N�E��u�e�d�d�g�m�F��H���T��
P��E��d�e�d�d�g�m�U���K���D��^�E��d�e�e�w�w�}�W��J���V��_�E��e�e�e�y�o�i�J���I����W��^�D��y�m�`�h�w�m�F��H����W��L����u�g�u�k�u�m�G��I����V��B��G���k�w�e�e�f�l�F��H���^��S�W��e�d�e�e�f�m�F��s���T��
P��E��d�d�d�e�f�m�U���J���D��^�D��e�e�d�w�w�n�W���[����V��_�E��w�u�u�u�o�o�J���I����V��_�D��y�m�f�h�w�m�F��I����V��L�M��h�u�e�d�g�l�G��H����FǻN��F���k�w�e�d�g�l�G��H���^��S�W��d�e�d�d�f�l�F��A���F�_�D��e�d�d�d�{�W�W���J���D��_�E��e�d�d�w�w�n�W���[����W��^�E��w�u�a�u�i��G��H����W��^��U���u�m�d�h�w�m�F��H����V��L�M��h�u�e�d�f�m�G��I����F��N��U��d�d�e�d�g�l�G���Y���^��S�W��d�e�d�e�g�l�F��A���F�_�E��d�e�e�e�{�e�A��Y����W��_�D��d�y�_�u�w�i�W���[����V��^�E��w�u�a�u�i��G��H����W��_��U��u�k�w�e�f�l�F��I����J�N��M��h�u�e�d�f�m�F��H����F��N��U��d�d�d�e�f�l�G���Y����X�^�D��e�e�e�d�u�}�W���A���F�_�D��d�e�d�e�{�e�C��Y����V��^�D��e�y�m�`�j�}�G��I����W��^�Y�ߊu�u�`�u�i��F��I����V��^��U���u�k�w�d�g�m�G��H����J�V��K���d�e�e�d�g�m�F��U���F��N��U��e�e�d�d�g�m�G���Y����X�_�E��e�d�d�d�u�}�A���G����V��_�D��e�w�u�u�w�e�E��Y����V��_�E��d�y�m�f�j�}�G��I����W��^�Y��a�h�u�e�g�m�F��I����D�=N��U��u�k�w�d�g�l�F��I����J�X��K���d�e�e�e�f�m�G��U����[�^�E��d�e�e�d�f�q�}���Y����X�_�D��d�d�e�e�u�}�A���G����V��^�E��e�w�u�b�w�c�U��I����W��^�W���u�u�m�d�j�}�G��H����V��_�Y��g�h�u�e�g�l�G��I����D�Y�H���e�e�d�e�f�l�G��[��ƹF� Z��K���d�e�d�d�g�m�G��U����[�^�E��e�e�e�e�f�q�O��D���V��_�D��e�e�y�_�w�}�@���G����V��_�E��d�w�u�b�w�c�U��I����W��^�W���b�u�k�w�f�l�G��I����V�d��U��e�h�u�e�g�m�G��H����D�V�H���e�e�e�e�f�m�F��[����F�L�E��d�e�d�d�g��W���Y����[�^�D��d�e�e�e�f�q�O��D���V��_�E��e�d�y�m�b�`�W��I����V��^�D���_�u�u�m�w�c�U��H����W��^�W���m�u�k�w�f�l�F��H����V�V�U��w�d�d�d�f�l�F��I���F�V�H���e�e�e�d�f�m�F��[����F�L�E��d�e�e�d�f��W��Y���W��_�D��e�e�w�u�w�}�O��D���V��^�D��e�d�y�m�d�`�W��I����W��^�E���m�a�h�u�g�m�F��I����V��NךU���l�u�k�w�f�l�G��H����V�V�U��w�d�d�e�g�m�G��I���
Q�	N��D��e�d�e�d�g�m�[�ԜY����F�L�E��d�d�e�d�g��W��Y���W��_�E��d�e�w�u�g�}�I���H����V��_�E���u�u�u�l�f�`�W��I����V��_�E���l�g�h�u�g�m�F��H����V��N�F��u�e�e�d�f�m�G��I���9F�W�U��w�d�d�d�g�l�F��H���S�	N��D��d�d�d�d�f�m�[��O���V��_�D��e�d�e�y�]�}�W��Y���W��^�E��d�e�w�u�g�}�I���H����V��^�E���u�e�u�k�u�l�G��H����W��B��U���l�e�h�u�g�l�G��H����V��N�D��u�e�d�e�f�m�F��H���
W��
P��E��e�d�d�d�g�l�U���Y���U�	N��D��e�d�d�d�g�l�[��M���V��^�D��e�d�d�y�n�h�J���I����V��_�D��y�_�u�u�f�}�I���H����V��^�E���u�d�u�k�u�l�G��H����W��B��D���k�w�d�e�f�l�F��H���l�N�L��u�e�d�e�f�m�G��H���
T��
P��E��e�d�d�e�g�m�U���K���D��^�D��e�e�d�w�w�}�W��K���V��^�D��d�d�d�y�n�n�J���I����V��_�E��y�l�a�h�w�m�F��I����V��L����u�g�u�k�u�l�G��H����V��B��G���k�w�d�e�g�l�G��H���_��S�W��e�e�d�d�f�l�F��s���
T��
P��E��d�d�e�d�f�l�U���K���D��^�D��e�d�e�w�w�n�W���[����V��_�D��w�u�u�u�n�l�J���I����W��_�E��y�l�g�h�w�m�F��I����V��L�L��h�u�e�d�f�m�F��H����FǻN��F���k�w�d�e�f�m�F��I���_��S�W��e�d�d�d�g�m�G��@���F�_�D��d�e�e�e�{�W�W���J���D��^�D��d�e�e�w�w�n�W���[����W��^�E��w�u�f�u�i��F��H����W��_��U���u�l�e�h�w�m�F��H����W��L�L��h�u�e�d�f�l�F��I����F��N��U��d�e�e�e�f�m�F���Y���_��S�W��d�e�e�e�g�m�F��@���F�_�E��d�e�e�d�{�d�B��Y����V��^�E��d�y�_�u�w�i�W���[����V��^�D��w�u�a�u�i��F��I����W��^��U��u�k�w�d�f�m�G��H����J�N��L��h�u�e�d�g�l�F��H����F��N��U��d�e�d�e�g�l�G���Y����X�_�E��e�e�d�d�u�}�W���@���F�_�E��e�d�d�e�{�d�D��Y����V��^�E��d�y�l�a�j�}�G��I����W��^�Y�ߊu�u�`�u�i��F��H����W��_��U���u�k�w�d�f�l�F��I����J�Y��K���d�d�d�d�f�l�F��U���F��N��U��d�e�e�d�f�m�F���Y����X�_�E��d�d�e�e�u�}�A���G����W��^�E��d�w�u�u�w�d�F��Y����V��_�E��e�y�l�g�j�}�G��I����V��^�Y��f�h�u�e�f�m�F��H����D�=N��U��u�k�w�d�f�l�F��I����J�[��K���d�d�d�d�g�l�F��U����[�^�D��d�d�d�e�f�q�}���Y����X�_�D��e�e�e�e�u�}�A���G����W��^�E��e�w�u�c�w�c�U��H����W��^�W���u�u�l�e�j�}�G��H����V��_�Y��d�h�u�e�f�l�G��I����D�Y�H���e�d�d�e�f�m�F��[��ƹF� ]��K���d�d�e�d�f�m�G��U����[�^�D��e�e�e�d�g�q�N��D���W��_�D��e�e�y�_�w�}�@���G����W��^�D��e�w�u�b�w�c�U��H����V��_�W���b�u�k�w�f�l�G��H����W�d��U��l�h�u�e�f�l�F��H����D�V�H���e�d�d�d�g�m�F��[����F�L�D��d�d�e�e�f��W���Y����[�^�D��d�d�e�d�g�q�N��D���W��_�D��e�d�y�l�c�`�W��H����V��_�E���_�u�u�m�w�c�U��H����W��^�W���m�u�k�w�f�l�F��I����W�W�U��w�d�d�d�g�m�F��H���F�V�H���e�d�d�e�f�l�G��[����
F�L�D��e�e�e�d�f��W��Y���W��_�E��d�d�w�u�w�}�N��D���W��^�D��e�d�y�l�e�`�W��H����W��_�E���l�f�h�u�g�l�F��H����V��NךU���l�u�k�w�f�l�F��H����V�W�U��w�d�d�d�f�l�F��H���
P�	N��D��d�e�e�d�f�m�[�ԜY����F�L�D��d�e�d�d�f��W��Y���W��_�E��e�e�w�u�n�}�I���H����V��_�D���u�u�u�d�g�}�I���H����V��_�E���u�e�d�h�w�m�F��H����W��L�D��u�k�w�d�f�l�G��H����J�N��D��u�k�w�d�f�l�G��H����J�^�H���e�d�d�d�g�m�F��[����S�	N��D��d�d�e�e�g�m�[�ԜY����P�	N��D��d�d�e�d�g�m�[��I���D��_�D��e�d�d�w�w�m�O��Y����W��^�E��e�y�_�u�w�m�N��Y����W��^�D��d�y�d�d�w�c�U��H����V��_�W���e�d�h�u�g�l�F��H����V��NךU���e�g�h�u�g�l�F��H����W��N�D���k�w�d�d�f�l�G��H���W��N��U��d�d�d�d�g�m�F���Y���W��N��U��d�d�d�d�g�l�F���Y����[�^�D��d�d�d�e�f�q�F��Y���W��_�D��e�d�w�u�w�}�F��Y���W��_�D��d�d�w�u�g�d�J���I����W��_�E��y�d�g�u�i��F��H����W��^��U���u�d�g�u�i��F��H����W��^��U��g�h�u�e�f�l�F��H����D�^�U���d�g�h�u�g�l�F��H����W��G���!�<� �0���!���7����t/��r<��0����u�u�!�>�:�}�����Ɠ9��X�����&�
� �'��g�������R��G�����;�u�u�u�6�9�G���	���R��UחX���!�0�<�u�%�3����&����F�N��U��
����u����P����V��^��D���=�;�u�u�w�}�W�������G��S�����'�u�k�r�p�f�W���YӃ��VFǻN��U���u�4�1�e�#�-�K�������9F�N�����3�_�x�,�#�8��������R��X �����'�6�&�n�]�8��������@9��V��D���'�6�&�u�6�9�F�������9F�N�����
�8�u�h�6�9�F�ԑT����[��DN�����4�0�:�3�w�}�WϷ�Yۥ��e9��c+��'´�1�d�u�u�2�����H�Ƹ�VǻN��U���u�4�1�d�#�-�K�������@F�I�\�ߊu�u�u�9�2�W�W���Y�����E_�����h�4�1�d�]�}�W����ƥ�l�D�����&�!�4�&�6�8�����Ƽ�\��DUװ���8�4�6�&�m�-����
�ί�XO�=�����u�u�<�u�4�6����Ӈ����S��D���!�0�_�u�w�}�W���Q����F�G�����_�u�u�u�w�}�W��E�ơ�^N��y8��;����}�1�'��0�^��s���F�R ����u�u�u�u�>�}���D����F��R ��U���u�u�u�u�&�}�Jϳ�ۥ��e9��c+��'´�1�d�!�%�~�}�W���Y����]��QUךU���;�u�3�_�9�}����
��ƓV��E�����<�'�'�u���}���Y������h�����d�a�4�9�]�8����Y����P��q��*���d�>�'�
�w�.�W�������Z�=N��U���u�4�4�<�#�}�W���<����	[�UךU���u�u�1�'�$�����Cӯ��v!��T��D��n�u�u�u�w�����
����[F��~ ��2���o�u�d�n�w�}����Y���F�N�����o��u����>��Y���F��[��U��������W�W���Y�ƭ�W��D^��U���������4���Q����V��^
��U���u����g�f�W���Y����VV�'��&������_�w�}�W���I����f2��c*��:���
�����)� ������"��y:��E��u�u�u�u�6�9����Y�ƅ�5��h"��<�������3�8�������F��` ��U���_�u�u�u�w�8�W���7ӵ��l*��~-�U���u�u�$�u�w��W���&����p9��t:��]���4�<�!�u�w�}�8���6���l��SN�����n�_�'�=�#�>��������\ ��\��C���3�e�3�d��<������F��Z�����8�g�e�f���(���H����A9��E���ߊu�u�u�u�8�)�_���Y���F���U���������}���Y���F�V
��E���u��
���(���-����F�N��U���6�e�o��w�	�(���0��ƹF�N��U���e�o�����;���:����g)��=N��U���u�u�u�1�%�}�W���*����|!��h8��!���_�u�u�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�w�}����Y����`2��{!��6�����|�_�w�}��������V��=dװ���;�u�u�8�e�m�Dۘ�&ù��W��V��G���8� �o�u�8�-����Y����P��q��*���d�>�'�
��2�}���Y������FךU���u�u�9�u�i�>��ԜY���F��S�H���1�'�&�e�]�}�W���Y����X��R^�U���u�u�$�u�i�,�[���Y�����E_��Kʴ�1�0�&�y�w�}�W������F��BךU���u�u�d�h�w�l�L����ƭ�P��R����_�