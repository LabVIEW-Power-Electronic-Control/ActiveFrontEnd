-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�M���� ^��1��@���
�
�e�
������
���F��Y���ߊu�u�u�u�w�}���� ���F��D�����h�w�9�6�u�}�W���Y���F��@�����u�o�<�!�0�/�M���K��ƹF�N��U���"�1�=�u�w�g�������F��d��U���u�u�u�8�:�.����Y����]��R��H��u�u�|�u�w�}����Y���F�N�����e�u�u�o�>�}��������E��X�����=�d�1�"�#�}�^���Y���F���U���u�u�u�;�$�9������ƹF�N��U��u�u�u�u�w�(�W���&����P9��T��]���1�=�d�1� �)�W���s���F�N����u�u�o�<�w�)�(�������P�������d�1�"�!�w�t�W���Y���F��R_��U���u�u�;�&�3�1����Y���F�N��D���u�u�u�u�9�.��������V��EF�����x�u�:�;�8�m�L�ԜY���F�@�U���u�o�<�u�#�����B���F�N�����u�u�u�u�w�3��������l�N�U��1�0�!�!�l�W�}�������G����U���8�a�c��o��(���&����lU��h��*���u�&�_�&�0�<�W���ù��CF��D�����6�#�6�:��*����Hӂ��]��G����0�8�8�4�%�$��������V��XN�����/�x�|�:�w�)�(�������P��F�����x�u�:�;�8�m�L���������^��ʧ�8�o�8�8�6�/���Yۉ��V��	F�����h�r�r�|�]�<��������J��V�����o�&�'�;�l�W��������@��E�����u�3�'�8�m�+�����ƥ�D��X�����n�4�!�<�"�8����
����\��C�����!�'�7�!�w�<�(����ƣ���T�����7�0�<�u�2�����s����Z��RN�� �����
���	�%���4����\��C���ߠ7�2�;�_�]�8��������@9��V��E���'�6�&�u�6�9�G�������9F�N�����
�8�u�h�6�9�G�ԑT����[��DN�����4�0�:�3�w�}�WϷ�Yۥ��e9��c+��'´�1�e�u�u�2�����H�Ƹ�VǻN��U���u�4�1�e�#�-�K�������@F�I�\�ߊu�u�u�9�2�W�W���Y�����E^�����h�4�1�e�]�}�W����ƥ�l�D�����&�!�4�&�6�8�����Ƽ�\��DUװ���8�'�
�6�2�.�G�������@F��[��U��2�;�_�u�w�;�_���^����GF��SN����r�r�u�=�9�}�W���Yӏ����S��D���!�0�u�u�w�}�W���Yӗ��[��V��:�������6�9�G���	����9F�N��U���u�3�_�u�w�3�W���s����C��R�����
�0�:�,�6�>����CӖ��P��F�����_�0�<�u�w�}��������E����U���u�u�d�|�#�8�}���Y���Z �T�H��r�u�=�;�]�}�W���Y���Z �@�H��r�u�=�;�]�}�W���Y���F�E��6���
�����9����Y����]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�3�_�9�}����
��Ɠ9����N�ߠ�7�4�,���L��ӯ��vH��S1�����d�c�{�9�l�W���� Ӌ��P��V��E���`�3�
�
�g��(���
�����R��U�ߊu�u�u�u�6�<����Y�ƅ�g#��eN�U��_�u�u�u�w�9����+����\��y:��0���h�a�_�u�w�}�W�������Z��T��;����u�h�g�l�}�WϮ����F�N�����!�o��u���8���B���F���U���������}���Y���R��R��U���������!���6�΍�W��D9�����u�u����m�L���Y�����T��;ʆ�����]�}�W���Y���)��=��*����
�����������W��x9��:��n�u�u�u�w�<����
����z(��c*��:���
�����9��������F��s!��!���|�_�u�u�w�}����Y����g"��x)��N���u�u�u�"�f�g�>���-����t/��=N��U���u�d�o��w�	�(���0����p2��*�����!�u�u�u���8��P���WF��C��N���'�=�!�6�"�8����Y����uR��/����3�`�3�
��m�(���Y��ƹF��X�����u��e�l�d�;�G���L����9��1��E���8�<�_�u�w�}�W�����ƹF�N��U���9�u�u����;���:���F�N��Uʴ�1�e�o��w�	�(���0����p2��d��U���u�u�u�6�g�g�>���-����t/��=N��U���u�u�u�e�m��#ύ�=����z%��r-��'�ߊu�u�u�u�w�}����Y�ƅ�5��h"��<������_�w�}�W���Y�Ư�F��~ ��!�����n�u�w�}�W���Yӂ��	F��=��*����
����W�W���Y���F��N�<����
���~�W�W����Ư�^��R ���ߠ7�2�;�u�w�0�C��8�ު�9��1��*ߊ�e�
�
�
�6��W�������]����E���f�3�e�3�b�;�(ځ�Iƹ��9��Zd��Uʥ�'�u�4�u�]�}�W���Y����X��[�U���u�u�4�1�g�`�W�������l�N��Uʶ�e�h�u�0�{�}�W���Yӗ��X��BךU���u�u�1�'�w�c��������9F�N��U���u�k�6�d�]�}�W���Y���F��d��U���u�"�d�h�w�8�^�Զ����A��C�� ���_�_