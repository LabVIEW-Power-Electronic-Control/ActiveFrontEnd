-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��b�d�l���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�4�0��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�^ �����
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W�������T��h��U���������!���6���F��@ ��U���_�u�u�;��3�������/��d:��9�������w�n�W������]ǻN�����;�0�b�0�c�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��a��R1�����o��u����>���<����N��
�����e�n�u�u�>�����&Ĺ��F��~ ��!�����
����_������\F��d��Uʼ�
�4�2�
���W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V �����!�:�
�g�2�m�Mϗ�Y����)��tUךU���;��;�4��3����H����F��~ ��!�����
����_������\F��d��Uʼ�
�4� �9�8�)����K����\��yN��1�����_�u�w�3�:�������G��h_����o��u����>���<����N��
�����e�n�u�u�>���������A	��\��*���u������4�ԜY�ƥ�l+��B�����:�
�g�0�b�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��~��V�����9�d�
�
�w�}�9ύ�=����z%��N�����4� �9�:�#�2�(������/��d:��9�������w�n�W������]ǻN�����<�&�a�0�g�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��t��D1����o��u����>���<����N��
�����e�n�u�u�>�����&ǹ��F��~ ��!�����
����_������\F��d��Uʼ�
�4�;�
���W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V��*ފ�
�u�u����;���:����g)��]����!�u�|�_�w�}��������l��T��;ʆ�������8���J�ƨ�D��^����u�;��<�$�i���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF��Y1�����a�0�b�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϷ�&����G9��N��U���
���n�w�}����/�ԓ�lV�'��&���������W��Y����G	�UךU���;��
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƥ�l6��1��G���u��
���(���-��� W��X����n�u�u�<���E���J����}F��s1��2������u�d�}�������9F���&���
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���*����V9��N��U���
���
��	�%���Hӂ��]��G�U���4�
�0� �9�m�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���R��R����o������0���/����aF�N�����u�|�_�u�w�-��������	F��cN��1��������}�D�������V�=N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӇ��A��E ��U��� �u��
���(���-��� W��X����n�u�u�4��8����L����f2��c*��:���
�����l��������l�N��*��� �;�c�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���	����F�� N�:���������4���Y����W	��C��\�ߊu�u�%�'�#�/�(���Y����`2��{!��6�����u�f�w�2����I��ƹF��G1�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}��������}F��s1��2���|�_�;�n�]�<��������VF��_�����e�c�`�d�1�m�����ƹF��X �����4�
�:�&��2����Y�Ɵ�w9��p'��O���d�n�u�u�4�3����Y����\��h�����u�u��
���W��^����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-�$�������^9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��1����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�e�d�g�f�W�������R��V��!���a�3�8�f�m��3���>����v%��eN��Bʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
��&�b�;���Cӵ��l*��~-��0����}�b�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6��#���O����lS�=��*����
����u�@Ϻ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������l��h��*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1��*���
�&�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�f�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'��(���I����l_�=��*����
����u�@Ϻ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������l��1����u�u��
���(���-��� Q��X����u�h�w�e�g�m�G��I����V��^�E��e�e�e�e�g��}���Y����G����&���!�g�3�8�f�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�f�m�G��I����l�N�����;�u�%���)�D�������	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W���*����R��D��F��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��_�E��e�e�e�e�l�}�WϽ�����GF��h=����
�&�
�a�m��3���>����v%��eN��Bʱ�"�!�u�|�m�}�G��I����V��^�E��e�d�e�e�g�m�G��I��ƹF��X �����4�
��&�f�����L����g"��x)��*�����}�b�3�*����P���V��^�E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����U��X��U���
���
��	�%���Nӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��h��M���8�d�u�u���8���&����|4�Y�����:�e�u�h�u�m�G��I����V��^�D��e�e�e�e�g�m�G���s���P	��C��U����
�!�l�1�0�F���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'��(���I����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��_�����e�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�g�
�&��l�Mύ�=����z%��r-��'���b�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
��.�E܁�
����\��c*��:���
�����j��������\�^�E��e�e�e�e�f�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����GT��Q��G���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1��*���`�3�8�g�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��_�E��e�e�e�e�g�m�G��I����F�T�����u�%��
�#�k����K����`2��{!��6�����u�f�w�2����I����D��^�E��e�d�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}����&����l ��h\�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��c1��GҊ�&�
�b�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
��&�g��.�(��Cӵ��l*��~-��0����}�b�1� �)�W���C���V��^�D��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6��#���Jù��^9��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��`2��C]�����f�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�g�3�:�n�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%����������F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��h��*��o������!���6���F��@ ��U���o�u�e�e�f�m�G��I����V��^�E��e�e�e�e�g�f�W�������R��V��!���f�
�&�
�c�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
��$�n�(���&���5��h"��<������}�`�9� ���Y���F�_�E��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)����-����9��Z1�U����
�����#���Q����\��XN�U��w�d�e�e�g�m�G��I����V��^�E��e�e�e�w�]�}�W���
������d:�����3�8�f�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�F��Cӵ��l*��~-��0����}�u�:�9�2�G���D����l�N�����;�u�%�6�9�)���&���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�rF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��_�W�ߊu�u�:�&�6�)��������_��h\�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��_�E��n�u�u�6�9�)����	����@��A]��G���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�D��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y�����e�o�����4���:����V��X����u�h�w�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�d�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�f��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�m�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�l�G���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��[��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�E���_�u�u�:�$�<�Ͽ�&����G9��\��M��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��e�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�e�w�_�w�}��������C9��Y����
��o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�e�l�}�WϽ�����GF��h�����#�g�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�g��}���Y����G�������!�9�f�
��g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�l�G��Y����\��V �����:�&�
�#�e�o�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�l�G��[���F��Y�����%�6�;�!�;�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��H���9F������!�4�
�:�$��܁�Y�Ɵ�w9��p'��#����u�g�1� �)�W���C���V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����F��d:��9�������w�l��������\�^�N���u�6�;�!�9�}��������EU��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�D��u�u�6�;�#�3�W�������l
��1�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�D��n�u�u�6�9�)����	����@��A]��4��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����\��h��G���o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�d�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�d�w�]�}�W���
������T�����f�
�f�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�f�f�W�������R��V�����
�#�g�g�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�d�g�m�U�ԜY�Ư�]��Y�����;�!�9�c��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#�c�l�Mύ�=����z%��r-��'���f�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�k�(���Y����)��t1��6���u�c�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�E��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��H���9F������!�4�
�:�$�����J����g"��x)��*�����}�f�3�*����P���V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������$�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����W��_�����u�:�&�4�#�<�(���
���� 9��N��1��������}�EϺ�����O�
N��E���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Kӂ��]��G��H���e�w�_�u�w�2����Ӈ��P	��C1��G��o������!���6�����Y��E���h�w�e�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�e�u�W�W�������]��G1�����9�m�e�o���;���:����g)��Y�����:�e�u�h�u�m�G��I��ƹF��X �����4�
�:�&��+�D��Cӵ��l*��~-��0����}�g�1� �)�W���C���V��^�E��e�e�e�e�g��}���Y����G�������!�9�d�
�g�m�Mύ�=����z%��r-��'���a�1�"�!�w�t�M���H����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��[��A��o������!���6���F��@ ��U���o�u�d�e�f�m�G��I���9F������!�4�
�:�$��ׁ�?����g"��x)��*�����}�u�8�3���Y���W��_�W�ߊu�u�:�&�6�)��������_��h[�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�l�(��Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�n�u�w�>�����ƭ�l��D�����a�e�o����0���/����aF�N�����u�|�o�u�g�m�F��I����V�=N��U���&�4�!�4��2�����֓�\��c*��:���
�����}�������	[�^�E��e�w�_�u�w�2����Ӈ��P	��C1��DҊ���u�u���8���&����|4�Y�����:�e�u�h�u�l�F��H����W��_�����u�:�&�4�#�<�(���
����^��rN�&���������W��Y����G	�N�U��e�e�e�e�f�l�F��[���F��Y�����%�6�;�!�;�l�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�e�w�_�w�}��������C9��Y����
��e�e�g�g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#�e�l�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�h�B��*����|!��h8��!���}�u�:�;�8�m�W��[����D��N�����!�;�u�%�4�3����L���5��h"��<������}�w�2����I����D��^�N���u�6�;�!�9�}��������ES��T��!�����
����_�������V�S��E��e�n�u�u�4�3����Y����\��h��*���u��
����2���+����W	��C��\��u�e�e�e�l�W�W���������t=�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�e�e�e�u�W�W�������F��Q�����1�;�u�u�#�4��ԜY�ƭ�G��B�����0�6�1�;�w�;����*����\��^	��ʼ�u�;�;�w�]�}�W�������C9��P1������&�d�3�:�m�Mύ�=����z%��N�����4�u�%�&�0�?���Y�Ǝ�|*��yUךU���<�;�9�3���Gځ�&ù��W��D^��U���
���
��	�%���Y����G	�UךU���<�;�9�3���Gځ�&ù��F��d:��9����_�u�u�>�3�ϸ�&����9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�?�D��L����l��E��D��������4���Y����\��XN�N���u�&�2�4�w�?�D��L����l��T��!�����n�u�w�.����Y����lU��h��*���u�u��
���L���Yӕ��]��Q��*��
�
�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������Q9��^�����4�1�0�&�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������Q9��^�����6�e�o����0���s���@��V�����f�`�0�d�&�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h]��Eߊ�
�
�1�'�$�l�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h]��Eߊ�
�
�0�u�w�	�(���0��ƹF��^	��ʳ�
�
�e�
������Y����)��tUךU���<�;�9�3���Gځ�&¹��\��c*��:���
�����l��������l�N�����u�7�f�f�b�8�E�������F��d:��9�������w�l��������l�N�����u�7�f�f�b�8�E���I����g"��x)��N���u�&�2�4�w�?�D��L����l��N��1��������}�D�������V�=N��U���;�9�3�
��m�(���&����V��T��!�����
����_�������V�=N��U���;�9�3�
��m�(���&����	F��s1��2���_�u�u�<�9�1����&����V9��@�Oʆ�����]�}�W�������Q9��^�����1�u�u����>���<����N��
�����e�n�u�u�$�:�����Փ�
S��V
�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����&����l��T��!�����n�u�w�.����Y����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�?�D��L����W��D_��U���
���
��	�%���Y����G	�UךU���<�;�9�3���N������5��h"��<��u�u�&�2�6�}����H����D��N��1�����_�u�w�4��������_��h
�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-����M�Փ�F��d:��9�������w�n�W������]ǻN�����9�'�2�d�b�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��*���$��
�!�d�;���Y�Ɵ�w9��p'�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������V��c1��G݊�&�
�c�o���;���:���F��P ��U���&�2�7�1�f�j�MϜ�6����l�N�����u�'�
� �f�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����a�c�o����0���/����aF�N�����u�|�_�u�w�4��������T9��R��!���g�
�&�
�d�g�$���5����l�N�����u�%�&�2�5�9�F��CӤ��#��d��Uʦ�2�4�u�!�d�l�Oׁ�I����g"��x)��*�����}�d�3�*����P���F��P ��U���
�a�g�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�f�
�&��o�Mύ�=����z%��N�����4�u�%�&�0�?���@����|)��v �U���&�2�4�u�'�.��������l��1����u�u��
���L���Yӕ��]��V�����1�
�l�u�w��;���B�����Y�����0�0�
�
�2�9����&����
V��N�&���������W������\F��d��Uʦ�2�4�u� ���Bց�����V��B1�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����J����l��E1����c�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ��Փ�P��V
��*���
� �a�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h]��@���4�1�
�0��n�@��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��[��*��m�4�1�
�2����O����	F��s1��2������u�f�9� ���Y����F�D�����!�f�d�m��9��������F��d:��9�������w�l��������l�N�����u� �
�
�o�i����&����U��Z��F��������4���Y����\��XN�N���u�&�2�4�w�(�(܁�A�ғ�W��E��G��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������U��N�&���������W������\F��d��Uʦ�2�4�u�
��8�(��L����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$���݁�
����	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������F9��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)��������F��d:��9�������w�k�W������]ǻN�����9�0�<�6�9�h����M�ѓ�F��d:��9�������w�m��������l�N�����u�'�
�:�2�)����Hƹ��9��h_�G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������G��h\�*���
�0�
�a�b�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����I����q)��r/�����u�<�;�9�2�4����M����R��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�����Jù��\��c*��:���
�����}�������9F������4�
�<�
�$�,�$����ԓ�@��N�&������_�w�}����Ӈ��@��U
��F��o�����W�W���������C��ي� �d�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��^	������
�!�f�1�0�F���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����l5��D�*���
�f�o����0���s���@��V�����2�7�1�f�d�g�5���<����F�D�����%�&�2�6�2��#���Hƹ��^9��T��!�����n�u�w�.����Y����Z��S
��C���u����l�}�Wϭ�����Z*��^1�����:�
�c�3��h�N���Y�Ɵ�w9��p'��#����u�g�1� �)�W���s���@��V��9���
�:�
�:�'�l�(���&����\��c*��:���
�����}�������9F������4�
�<�
�$�,�$����ѓ�@��N�&������_�w�}����Ӈ��@��U
��F��o�����W�W���������h]�����`�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��*��d�o�����4���:����P��S�����|�_�u�u�>�3�ϻ�����WT��B1�Aي�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����
9��T��!�����
����_������\F��d��Uʦ�2�4�u�%�$�:����&����GW��Q��D���u��
���f�W���
����_F��h��*���
�e�u�u���6��Y����Z��[N�����d�c�
�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�g�
�$��N��*����|!��d��Uʦ�2�4�u�%�$�:����M���$��{+��N���u�&�2�4�w����� ����S��R	��@��o������!���6���F��@ ��U���_�u�u�<�9�1����J���� 9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�-��������`2��C\�����g�u�u����>��Y����Z��[N��*���
�1�
�f�w�}�8���8��ƹF��^	��ʴ�
�<�
�&�&��(���K����lT��N��1�����_�u�w�4��������T9��S1�D������]�}�W�������F ��hW�*���
�e�o����0���/����aF�N�����u�|�_�u�w�4��������l ��h"����
�
�
�0��h�A��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��������;� �
�c�o����N�Փ� F��d:��9�������w�n�W������]ǻN�����9�3�
���o�8���Aǹ��A��[�U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������Q��N�&���������W������\F��d��Uʦ�2�4�u�8��o����K����	F��s1��2������u�g�9� ���Y����F�D����� �
�
�f�d�8�G���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����!��'��8��F���I����lT��N�&���������W��Y����G	�UךU���<�;�9�4��4�(�������@��h��*��o������}���Y����R
��G1�����1�a�l�o���2���s���@��V�����2�6�0�
��.�Eف�
����\��c*��:���n�u�u�&�0�<�W���
����W��W��U�����n�u�w�.����Y���� 9��_��*ڊ�e�o�����4���:����V��X����n�u�u�&�0�<�W�������A9��X��@���e�'�2�g�g�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������D�����
��&�g��.�(��Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������B9��h��E���8�g�u�u���8���B�����Y�����<�
�1�
�n�}�W���5����9F������3�
����(�(�������U��N�&���������W��Y����G	�UךU���<�;�9�3���2�������l��h\�C��������4���Y����W	��C��\�ߊu�u�<�;�;�?����H����V9��F^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�;�1�(���&����lT��R1�����g�f�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z��D��&���!�d�3�8�d�}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�7�1�n�F��&����BV�=��*����
����u�FϺ�����O��N�����4�u�9�9��2�(���	����V9��E��G��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ғ�F9��[��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������S��N��1��������}�GϺ�����O��N�����4�u�8�
�g�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����8�
�e�'�0�o�B���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
�
� �f�j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�d�<�'�0�o�A���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
�
� �e�m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�e�<�'�0�o�A���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
�
� �e�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�l�<�'�0�o�@���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���f�
�
� �e�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�b�<�'�0�o�@���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����F��a�
�
�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������~ ��-���!�'�
�a���(���&����\��c*��:���
�����l��������l�N�����u�!�f�d�c��(ށ�I����g"��x)��*�����}�d�3�*����P���F��P ��U�������#�/�(��&����A��Y�U����
�����#���Q����\��XN�N���u�&�2�4�w�)�D��MŹ��9��T��!�����
����_������\F��d��Uʦ�2�4�u�9���/�������S��R1�����g�e�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����lW��1��D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���0����r4��R��D���0�d�'�2�e�l�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��[��*��m�$�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����}"��v<�����b�
�0�
�`�h�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��[1��1����!�'�
�b��(߁�����V�=��*����
����u�FϺ�����O��N�����4�u�9����%�������9��1����a�u�u����>���<����N��
�����e�n�u�u�$�:��������v>��e����a�0�e�'�0�o�B���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*������0�:�l�C���H����lT��N�&���������W��Y����G	�UךU���<�;�9�<�d�;�(��N����	F��s1��2������u�e�9� ���Y����F�D�����
�
�0�
�`�n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��*���$��
�!�b�;���Y�Ɵ�w9��p'�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1����Jǹ��lT��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������P��N��1��������}�A�������V�=N��U���;�9�0�<�4�3�F���&����l��N��1��������}�GϺ�����O��N�����4�u�
�
�"�o�Cف�K����g"��x)��*�����}�u�8�3���B�����Y�����'�2�g�l�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�f�
�$��A��*����|!��d��Uʦ�2�4�u�%�$�:����L���$��{+��N���u�&�2�4�w�0�(�������T��N�&���������W��Y����G	�UךU���<�;�9�!�'�n�(���&����\��c*��:���
�����n��������l�N�����u�-�!�:�3�;�(��I����	F��s1��2������u�g�9� ���Y����F�D����� �
�
�e���(�������\��c*��:���
�����}�������9F������7�3�f�f�b�8�G���I����g"��x)��N���u�&�2�4�w�(�(܁�Iƹ��9��T��!�����
����_������\F��d��Uʦ�2�4�u� ���Gځ�&ù��W��D_��U���
���
��	�%���Y����G	�UךU���<�;�9�7�1�n�D����֓�VW�=��*����n�u�u�$�:�������� V��R1����o������}���Y����R
��B��*��
�
�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������F ��h]�*���
�d�o����0���/����aF�N�����u�|�_�u�w�4��������lU��h��*���'�&�e�o���;���:����g)��_�����:�e�n�u�w�.����Y���� 9��1��D���e�o�����4�ԜY�ƿ�T����*ي�e�
�
�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h]��Eߊ�
�
�1�'�$�l�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Q1��F���0�d�6�d�m��3���>����F�D����� �
�
�e���(���Y�Ɵ�w9��p'�����u�<�;�9�5�;�D��L����l��N��1��������}�D�������V�=N��U���;�9�7�3�d�n�B���H����	F��s1��2������u�d�}�������9F������7�3�f�f�b�8�E�������F��d:��9�������w�l��������l�N�����u� �
�
�g��(݁�����`2��{!��6�ߊu�u�<�;�;�?����J�ӓ�lT��N�&���������W��Y����G	�UךU���<�;�9�7�1�n�D����ԓ�W��D�Oʆ�������8���Hӂ��]��G�U���&�2�4�u�"��(��&����P��N��1�����_�u�w�4��������lU��h��*���u�u��
���L���Yӕ��]��U��F��`�0�g�1�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Q��1�@���g�$�u�u���8���&����|4�_�����:�e�n�u�w�.����Y���� 9��1�����&�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ��Փ�_��R^��U���
���n�w�}�����Ʈ�U9��[�����0�&�u�u���8���&����|4�N�����u�|�_�u�w�4��������l_��h��U����
���l�}�Wϭ�����Q��1�L���d�o�����4�ԜY�ƿ�T����*ي�`�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӄ��lU��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;�?����H����R��R��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�;�D��Oʹ��F��d:��9����_�u�u�>�3�ϼ��Փ�P��V
�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����J����
9��N�&������_�w�}����ӄ��lU��X����o������}���Y����R
��B��*���l�1�u�u���8���&����|4�_�����:�e�n�u�w�.����Y���� 9��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;�?����K����V9��V
�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����J����9��1��E�������W�W���������h]��L���0�e�4�1�2�.�W���-����t/��a+��:���d�1�"�!�w�t�}���Y����R
��B��*��d�0�e�6�f�g�$���5����l�N�����u� �
�
�n�l�������5��h"��<��u�u�&�2�6�}����&����l��h
�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�"��(��H����l��N��1��������}�GϺ�����O��N�����4�u� �
��d�F���H����A��N�&���������W������\F��d��Uʦ�2�4�u� ���N����ד�VV�=��*����n�u�u�$�:��������_��h��*��o������!���6���F��@ ��U���_�u�u�<�9�1����J����9��1�����&�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ��Փ�
U��R1����o������}���Y����R
��B��*��d�0�d�"�f�g�$���5����l�N�����u� �
�
�n�l��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʷ�3�f�g�f���(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�� ���
�c�e�0�g�<����
����`2��{!��6�����u�d�3�*����P���F��P ��U���
�
�c�e�2�m���Cӵ��l*��~-�U���&�2�4�u�"��(��I����l��E��D��������4���Y����\��XN�N���u�&�2�4�w�(�(܁�O�֓�lV��R_��U���
���n�w�}�����Ʈ�U9��X�*���
�0�u�u���8���B�����Y�����f�d�g�
���F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*ي�c�e�0�e�&�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��Q1��D��
�
�
�1�%�.�G��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U��F��g�
�
�
�2�}�W���&����p]ǻN�����9�7�3�f�f�o�(���&����V��T��!�����
����_�������V�=N��U���;�9�7�3�d�l�E߁�&¹��F��d:��9����_�u�u�>�3�ϼ��Փ�T��R1����o������}���Y����R
��B��*��e�0�d�1�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Q��1�Gڊ�
�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӄ��lU��^��*ڊ�1�'�&�e�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�U9��_�����6�e�o����0���s���@��V�� ���
�d�
�
��m�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��B��*��
�
�
�1�%�.�F��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U��F��e�0�e�6�f�g�$���5����l�N�����u� �
�
�f��(߁�����`2��{!��6�ߊu�u�<�;�;�?����@�֓�lV��N�&���������W��Y����G	�UךU���<�;�9�7�1�n�N����֓�F��d:��9�������w�n�W������]ǻN�����9�7�3�f�n�m��������@��N��1��������}�FϺ�����O��N�����4�u� �
��l�(���&����	F��s1��2���_�u�u�<�9�1����J����l��h�����d�o�����4���:����W��X����n�u�u�&�0�<�W���&����9��1��D�������W�W���������h]��Dڊ�
�
�0�u�w�	�(���0��ƹF��^	��ʷ�3�f�l�e�2�l����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����l�e�0�d�&�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��Q1��D��
�
�
�1�%�.�G��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U��F��f�
�
�
�2�}�W���&����p]ǻN�����9�7�3�f�f�n�(���&����V��T��!�����
����_�������V�=N��U���;�9�7�3�d�l�D܁�&ù��F��d:��9����_�u�u�>�3�ϼ��Փ� U��R1����o������}���Y����R
��B��*��f�0�e�1�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Q��1�Fي�
�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӄ��lU��]�����4�1�0�&�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������F ��h_�F���d�6�e�o���;���:���F��P ��U���
�
�f�f�2�l��������	F��s1��2������u�f�9� ���Y����F�D����� �
�
�f�d�8�F���H����g"��x)��N���u�&�2�4�w�(�(܁�J�Փ�lW��R_��U���
���n�w�}�����Ʈ�U9��]�*���
�d�o����0���/����aF�N�����u�|�_�u�w�4��������lW��1��D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���J����9��S�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�1�(܁�O�ޓ�VV�=��*����n�u�u�$�:�����Փ�^��V
�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����&����l��T��!�����n�u�w�.����Y����lW��1��D�������W�W�������
��1�MҊ�d�o�����4���:����U��S�����|�_�u�u�>�3�ϲ�&����P��h^�����&�e�o����0���/����aF�
�����e�n�u�u�$�:�����Փ�R��R1����o������}���Y����R
��C1��D��
�
�
�1�%�.�F��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��[��*��c�0�e�6�f�g�$���5����l�N�����u�!�f�d�c��(߁�����`2��{!��6�ߊu�u�<�;�;�1�(܁�A�Г�lV��N�&���������W��Y����G	�UךU���<�;�9�9���O����ד�W��D�Oʆ�������8���Hӂ��]��G�U���&�2�4�u�#�n�F��&����P��N��1�����_�u�w�4��������^��h��*���'�&�d�o���;���:����g)��_�����:�e�n�u�w�.����Y����lW��1��D���d�o�����4�ԜY�ƿ�T����F��a�
�
�
�2�}�W���&����p]ǻN�����9�9�
�
�o�k��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʹ�
�
�c�`�2�m��������	F��s1��2������u�f�9� ���Y����F�D�����!�f�`�l���(���Y�Ɵ�w9��p'�����u�<�;�9�;��(��L����l��N��1��������}�D�������V�=N��U���;�9�9�
��k�B���I����A��N�&���������W������\F��d��Uʦ�2�4�u�!�d�h�Nځ�&ù��F��d:��9����_�u�u�>�3�ϲ�&����
S��h^�����u��
���f�W���
����_F��h]��C���0�e�1�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ơ�lU��W�����$�u�u����>���<����N��
�����e�n�u�u�$�:�����Փ�_��R1�����0�&�u�u���8���&����|4�N�����u�|�_�u�w�4��������P��h��*���u�u��
���L���Yӕ��]��[��*��`�0�d�$�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����_��h[�@���d�4�1�0�$�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������
��1�Lߊ�
�
�0�u�w�	�(���0��ƹF��^	��ʹ�
�
�c�`�2�l� ��Cӵ��l*��~-�U���&�2�4�u�#�n�B��&����WW�=��*����
����u�FϺ�����O��N�����4�u�!�f�b�d�(���&���5��h"��<������}�f�9� ���Y����F�D�����!�f�`�l���(�������\��c*��:���
�����}�������9F������9�
�
�c�b�8�E���I����g"��x)��N���u�&�2�4�w�)�D��@ƹ��9��T��!�����
����_������\F��d��Uʦ�2�4�u�!�d�h�Nځ�&����W��D_��U���
���
��	�%���Y����G	�UךU���<�;�9�9���A����ԓ�VW�=��*����n�u�u�$�:�����Փ�_��R1����o������}���Y����R
��C1��@��
�
�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������G9��X�*���
�d�o����0���/����aF�N�����u�|�_�u�w�4��������lW��1�����&�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ��Փ�^��T�Oʆ�����]�}�W�������F ��h_�A���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����R��S
����o������!���6�����Y��E��u�u�&�2�6�}����&����l��T��!�����n�u�w�.����Y���� 9��Z�����u��
���f�W���
����_F��Q1��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����J���5��h"��<������}�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��\�Oʗ����_�w�}����Ӈ��l��R1�����d�
�
�0��n�A��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������
F��u!��0���_�u�u�<�9�1��������V��c1��M���8�b�o����0���s���@��V�����2�7�1�m�`�g�5���<����F�D�����d�'�2�d�`�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������D�����
��&�d��.�(��Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}�;���&����	��h�����f�l�o����0���/����aF�
�����e�n�u�u�$�:����	����l��F1��*���c�3�8�d�w�}�#���6����9F������4�
�<�
�3��@���Y����v'��=N��U���;�9�4�
�>�����*���� T��D��D�������W�W���������D�����m�m�o����9�ԜY�ƿ�T�������d�e�u�u���8���&����|4�N�����u�|�_�u�w�4��������T9��R��!���f�
�&�
�b�g�$���5����l�N�����u�%�&�2�5�9�O��CӤ��#��d��Uʦ�2�4�u�f�%�:�F��Y�Ɵ�w9��p'��#����u�d�1� �)�W���s���@��V�����2�6�0�
��.�Dׁ�
����\��c*��:���n�u�u�&�0�<�W���
����W��V��U�����n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��F���Y����v'��=N��U���;�9�4�
�>�����*����9��Z1�Oʆ�����]�}�W�������C9��P1����`�o�����}���Y����R
��Z��*���d�e�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������^��1��*���l�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��C���Y����v'��=N��U���;�9�4�
�>�����*����V��D��U����
���l�}�Wϭ�����R��^	�����c�u�u����L���Yӕ��]��C��Fڊ� �d�f�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������D�����
��&�g��.�(��Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}����7����V��V��*؊� �g�d�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��D��
�e�o����0���/����aF�N�����u�|�_�u�w�4��������F9��]��D��������4���Y����W	��C��\�ߊu�u�<�;�;�:����&����l��N��1��������}�D�������V�=N��U���;�9�2�%�1��C���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�
�a�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����a�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��D��
�e�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�G���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ӓ�F9��Y��E��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����R��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:��N���&����l��N��1��������}�D�������V�=N��U���;�9�!�%�`����L����\��c*��:���
�����l��������l�N�����u�8�
�m�1��B���	����`2��{!��6�����u�d�3�*����P���F��P ��U��� ����#�/�(�������W��N�&���������W��Y����G	�UךU���<�;�9�9�4�����L�ӓ�F��d:��9�������w�j��������l�N�����u�:�
�
�e�;�(��L����	F��s1��2������u�e�}�������9F������!�%�<�<�>�n�(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�<�>�4����L�ߓ�F��d:��9�������w�m��������l�N�����u�0�
�
�����@¹��\��c*��:���
�����i��������l�N�����u�8�
�f���(�������
9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(�������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(�������9��T��!�����
����_�������V�=N��U���;�9�'�!�e�4��������P��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	����F
��D1��*��d�%�u�u���8���&����|4�Y�����:�e�n�u�w�.����Y����~3�� ����
�;�0�%��o����O�ߓ�F��d:��9�������w�l�W������]ǻN�����9�!�%�<�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�d�
�
�"�l�Aށ�K����g"��x)��*�����}�u�8�3���B�����Y�����`�
� �d�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Cڊ� �d�m�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��[�� ��m�
�d�o���;���:����g)��Y�����:�e�n�u�w�.����Y����W��B1�Lي�f�o�����4���:����Q��X����n�u�u�&�0�<�W���H�ד�l��B1�Bي�f�o�����4���:����T��S�����|�_�u�u�>�3�Ϫ�	����Z9��h_�D���u�u��
���(���-��� V��X����n�u�u�&�0�<�W�������lQ��Q��B���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����2��x��Mފ�;�3��%��(�F��&���5��h"��<������}�c�9� ���Y����F�D�����0�
�8�c�>�;�(��L����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�b�>�;�(��H����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�m�>�;�(��N����	F��s1��2������u�g�9� ���Y����F�D������-� ��9�(�(�������W��N�&���������W��Y����G	�UךU���<�;�9�;�#�5�(���H����CT�=��*����
����u�W������]ǻN�����9�%��9��h����N�֓�F��d:��9�������w�n�W������]ǻN�����9�9�6��f����N����\��c*��:���
�����}�������9F������9�6��d��(�F��&���5��h"��<������}�e�9� ���Y����F�D�����8�
�
�g�>�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����8�
�
�f�>�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����
�4�g�b��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����:�
�
�`�1��O���	����`2��{!��6�����u�b�3�*����P���F��P ��U���
�
�c�3��e�N���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����<�<�
�
�d�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����8�
�
�a�>�;�(��@����	F��s1��2������u�g�9� ���Y����F�D�����
�4�g�b��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����:�
�
�b�1��O���	����`2��{!��6�����u�b�3�*����P���F��P ��U���
�
�m�3��e�B���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����<�<�
�
�c�;�(��@����	F��s1��2������u�g�9� ���Y����F�D�����8�
�
�`�>�;�(��L����	F��s1��2������u�g�9� ���Y����F�D�����:�'�&�
�"�l�O܁�K����g"��x)��*�����}�u�8�3���B�����Y�����=�`�3�
�o�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�� �����
� �d�e��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��C��C���
�m�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��h_�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����OĹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�0�-����M�Г�F��d:��9�������w�m��������l�N�����u�:�'�&��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʻ�!�=�b�3��d�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����e�3�
�l�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��D���
�l�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��h_�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Nʹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�F�������T��^1��*��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������_��R�����<�3�
�m�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z�����l�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lW��h
�����;�<�3�
�`�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�l�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��DҊ�
�0�:�2�9�;�(��L����	F��s1��2������u�g�9� ���Y����F�D�����8�
�f�3��d�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�
�
�"�l�Nށ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�l�<�1��N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�d�
��2�(���K����CT�=��*����
����u�W������]ǻN�����9�!�%�b��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�m�>�;�(��L����	F��s1��2������u�g�9� ���Y����F�D�����8�
�a�3��m�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����m�3�
�e�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��d1��9����!�d�c�1��G���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�<�8�
�
�"�o�A݁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�d�
��(�E��&���5��h"��<������}�f�9� ���Y����F�D�����0�
�8�g�����Nǹ��\��c*��:���
�����l��������l�N�����u�0�
�8�d��(���K����CU�=��*����
����u�FϺ�����O��N�����4�u��!�%�l�F���M����V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�1�����&���� 9��h\�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����9��Q��E���%�u�u����>���<����N��
�����e�n�u�u�$�:��������CS��^1��*��e�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G��1�����d�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��h_�F���6�1�u�u���8���&����|4�N�����u�|�_�u�w�4��������F9��]���������W�W���������D�����
��&�d��.�(��Cӵ��l*��~-�U���&�2�4�u�'�.��������
F��u!��0���_�u�u�<�9�1�������� P��G����������4���Y����\��XN�N���u�&�2�4�w�0�(�������T��G����������4���Y����\��XN�N���u�&�2�4�w�0�(�������Q��G����������4���Y����\��XN�N���u�&�2�4�w�0�(�������T��G����������4���Y����\��XN�N���u�&�2�4�w�-�9���
����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�
�<�
�1��e�N��;����r(��N�����4�u�%�&�0�?���@����q)��r/�����u�<�;�9�6���������T�,��9���n�u�u�&�0�<�W���
����W��X��U�����n�_�w�}��������^V�� [�L���
�4�1�&�5�n����K����9��Q��*���u��u�u�0�3����Q���F�'��Oʜ����_�w�}�W���,����r!��N��!����_�u�u�w�}����.����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�:�#�
�3���Cӯ��v!��G�U���%�'�u�_�w�}�W�������z(��c*��:���n�u�u�u�w�/����Cӯ��`2��{!��6�ߊu�u�u�u�>�m�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y���F��^ �Oʜ�u��
����2���+������Y��E��u�u�u�u�8�>����Y����g"��x)��*�����}�u�8�3���B���F���Oʜ�u��
���f�W���Y����\��N��!ʆ�������8���J�ƨ�D��^��\�ߊu�u�;�u�8�-����B��ƹF��X�����u�e�c�`�f�;�G�������]�� ��F؊�
�4�
�&�w��W�������Z�=N��U���u��o����%�ԜY���F��z1��4���o�����W�W���Y�ƨ�]V��~*��U������n�w�}�W�������d/��N�<�����_�u�w�}�W�������g.�'��0���u�n�u�u�'�/�W�ԜY���F��Y^��U���������4���Y����W	��C��\�ߊu�u�u�u�>�l�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y���F��X��Oʚ�������!���6���F��@ ��U���|�_�u�u�9�}��������9lǻN�����;�;�u�e�a�h�Fָ�I����C9��Y��G���d�d��_�w�}�������F�N��<���u����l�}�W���YӨ��l5��p+��U�����n�u�w�}�WϺ�ù��w2��N��!����_�u�u�w�}����.����\��y:��0��u�u�u�u�3�(�(���-����z(��p+��\�ߊu�u�:�!��}�W���Yӂ��F��~ ��!�����
����_������\F��d��U���u�1�;�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƣ�P	��T��;ʆ�������8���Mӂ��]��G�U���u�u�1� �w�}�"���-����t/��a+��:���e�1�"�!�w�t�^�ԜY�Ʃ�WF��Z�����_�_�u�u�8�-����Y�֍�S����*���
�7�f�f�b�8�Gϗ�s���T��E��]���u�u�u��#�
����Cӯ��v!��d��U���u��1�0�$�<����Y����t#��=N��U���u�1�'�&� �9���0����v4�d��Uʥ�'�u�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�%�.���0�Ɵ�w9��p'�����u�u�u�1�%�.�G��0�Ɵ�w9��p'��#����u�d�1� �)�W���s���F�T�Oʜ�u��
���f�W���Y����F��x;��&���������W��Y����G	�UךU���u�u�1�'�$�l�Mϗ�Y����)��t1��6���u�d�1�"�#�}�^�ԜY���F��N�<����
���l�}�W���Yӑ��\��yN��1�����_�u�w�}�W��Cӯ��`2��{!��6�����u�f�w�2����I���9F���U���%�;�;�n�]�}�WϽ�����]��/�@��3�e�3�f�1��(��Jӯ��F�P�����}�u�u�u�w��������/��r)��N���u�u�u��3�8��������z(��p+�����u�u�u�1�%�.� �������}2��r<��N���u�%�'�u�]�}�W���Y����	F��=��*����n�u�u�w�}��������}F��s1��2���_�u�u�u�w�9����I����}F��s1��2������u�g�9� ���Y����F�N����o��u����>��Y���F��N�:���������4���Y����W	��C��\�ߊu�u�u�u�3�/���Cӯ��`2��{!��6�����u�e�3�*����P���F�N��D���u��
���L���Y�����T��;ʆ�����]�}�W���Y���/��d:��9�������w�n�W������F�=N��U���u�:�%�;�9�f�}���YӅ��C	��Y��E��`�d�3�e�1�n����J����l��'��U���2�;�'�6��}�W���YӢ��R1��C��U�����n�u�w�}�Wϟ�����a��RN�<�����_�u�w�}�W�������Z��T��;����u�n�u�w�-����s���F�T��Oʜ�u��
���f�W���Y����V��T��;ʆ�����]�}�W���Y����V��T��;ʆ�������8���Hӂ��]��G�U���u�u�6�e�m��W���&����p]ǻN��U���e�o�����;���:����g)��]����!�u�|�_�w�}�W�������@W�'��&���������W������\F��d��U���u�6�d�o��}�#���6����9F�N��U���u�u�����0���s���F�S_��U���������4���Y����W	��C��\�ߊu�u�u�u�f�g�8���*����|!��h8��!���}�d�1�"�#�}�^���s���V��T�����!�_�_�u�w�2�����ơ�rP��_��*ڊ�
�
� �
��d�F���Iӯ��F�P�����}�u�u�u�w��������/��r)��N���u�u�u��3�8��������z(��p+�����u�u�u�1�%�.� �������}2��r<��N���u�%�'�u�]�}�W���Y����	F��=��*����n�u�u�w�}��������}F��s1��2���_�u�u�u�w�9����I����}F��s1��2������u�f�9� ���Y����F�N����o��u����>��Y���F��N�:���������4���Y����\��XN�N���u�u�u�4�3�8����Y����g"��x)��*�����}�u�8�3���B���F���U���������}���Y���D��N��U���
���n�w�}�W�������z(��c*��:���
�����}�������9F�N��U��o������0���/����aF�
�����e�u�n�u�w�8�Ͻ�����]��=d��Uʶ�8�:�0�!�:��@��@����U9��U��F��m�u��u�w�:������ƹF�N�����<�!�u�u���2��Y���F��S
�����;�0�o����%�ԜY���F��S�����!�u�u����W��Y����\��d��U���u�6�>�o��}�#���6����9F�N��U���0�u�u����;���:���F�N�����&�u�u����;���:����g)��^�����:�e�n�u�w�}�WϽ�I����}F��s1��2���_�u�u�u�w�m�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���F�V
�����u�u�����0���/����aF�
�����e�n�u�u�w�}���Cӯ��`2��{!��6�ߊu�u�u�u�2�}�W���*����|!��d��U���u�1�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y���)��=��*����
����u�FϺ�����O�d��Uʰ�1�6�8�:�2�)�}�Զ����9F���F��`�0�e� �m�>��������'��_����3�f�3�
��m�(���s���T��E�����}�u�u�u�w��������F��d��U���u��1�0�$�<����G����F�N��4���0�&�<�!�w�c�E�ԜY�Ƽ�A��V�����u�u�u�9�w�c������ƹF�N�����u�k�4�
�$�q�W���Y����W��D�H���7�f�f�`�2�m��������9F�N��U���u�k�3�
��m�(���&����9F�N��U��h�u�7�f�d�h������ƹF�N�����&�d�h�u�5�n�D����֓�W��D����u�u�u�0�w�c����&����V9��T����u�u�u�0�w�c����&����V9��@����u�u�u�d�j�}����J�ӓ�lV��G����u�7�f�f�b�8�F���CӅ��C	��Y��E��`�d�3�e�1�n����&����V9��N�����'�6�8�%��}�W���YӢ��R1��C��K��y�u�u�u�w�����
����VF�Z�U���u�u��1�2�.����Y���l�N�����4�u�_�u�w�}�W���Y����C9��\BךU���u�u�0�0�w�c����
��ƹF�N�����&�e�h�u�5�n�D����ד�W��D����u�u�u�0�w�c����&����V9��T����u�u�u�e�j�}����J�ӓ�lW��BךU���u�u�1�'�$�l�J����Փ�S��h_�����&�d�_�u�w�}�W���Y����Q9��^�����6�d�_�u�w�}�W���Y����Q9��^�����"�d�_�u�w�}�W��D�ƪ�lU��[��*ۊ�d�n�_�u�w�?�D��L����l3������;�u�e�c�b�l�����Փ�Q9��^����u�u�2�;�%�>����Q���F�*�����!�u�k�f�{�}�W���Yӧ��A��e����u�y�u�u�w�}�6�������W��
P��\���u�%�'�u�6�}�}���Y���P
��
P�����>�_�u�u�w�}����Y����C9��CBךU���u�u�1�'�$�m�J����Փ�S��h\�����&�e�_�u�w�}�W���Y����Q9��^�����6�e�_�u�w�}�W��D�ƪ�lU��[��*؊�e�_�u�u�w�}����
���F��h]��Eߊ�
�
�1�'�$�l�}���Y���P��
P�����f�`�0�g�4�l�}���Y���D��
P�����f�`�0�g� �l�}���Y���WW�	N��*ي�e�
�
�
�f�f�}���Y����lW��1��Oʶ�8�:�0�!�:��@��@����U9��Q��*��f�u�u�2�9�/�ϳ�	��ƹF�N�����<�!�u�k�d�q�W���Y����W��D�����h�u�y�u�w�}�Wϟ�����d��_N��U���u�u�%�'�w�<�W�ԜY���F��\N��U���6�>�_�u�w�}�W��������E�����u�u�u�1�%�.�G��Y����lW��1�����&�y�u�u�w�}���D�ƪ�lU��[����_�u�u�u�w�m�J����Փ�
S��F^�U���u�u�4�1�2�.�W�������_��h�����d�_�u�u�w�}����GӀ�� 9��]�����u�u�u�u� �l�J����Փ�
S��@����u�u�u�d�j�}����H����WW�=d��Uʷ�3�f�f�`�2�m�"������]����C���d�3�e�3�d�?����J�ӓ�lVǻN�����<�u�4�u�]�}�W���Y����d��_N��U��_�u�u�u�w�9����+����[�BךU���u�u�1�'�$�
����D����9F���ʸ�%�}�u�u�w�}����D�ƭ�l��d��U���u�'�&�!�j�}�������F�N�����&�u�k�7�1�n�D����֓�W��D����u�u�u�0�w�c����J����l��h��Y���u�u�u�$�w�c����J����l��h����u�u�u�1�%�.�F��Y���� 9��1��E���1�0�&�y�w�}�W������F��Q1��F���0�e�6�d�]�}�W���Y����X��B��*��
�
�
�0�{�}�W���Yӂ��X��B��*��
�
�
�d�]�}�W���Y���F��Q1��F���0�e�$�|�]�}�Wϼ��Փ�S��h_��U���:�%�;�;�w�m�A��Hʀ��l ��h��*ي�e�
�
�_�w�}�����ơ�CF�N��U����!��1�?�`�W��s���F�v
�����4�2�u�k�c�W�W���Y�ƍ�W��D9�����k�g�_�u�w�2�ϳ�	��ƹF�N�����k�4�
�9�{�}�W���YӔ��V�	N��*���y�u�u�u�w�<����
�����h]��Eߊ�
�
�1�'�$�m�}���Y���P��
P�� ���
�e�
�
��8�[���Y�����
P�� ���
�e�
�
��m�}���Y���R��R��U��7�3�f�f�b�8�F�������JǻN��U���0�u�k�7�1�n�D����ד�VW�N��U���"�d�h�u�"��(��&����D��=N��U���u�d�h�u�"��(��&����WW�N��U���$�u�k�7�1�n�D����ד�O��=N��U���
�
�e�
���W�������V��Z^��B��l�
�
�
��(�(܁�Iƹ��l�N�����6�8�%�}�w�}�W���=����Z��S�F���u�u�u�u��9��������X�d��U���u��1�0�$�4����G���F�G��U���u�_�u�u�w�}����GӇ��P
��=N��U���u�0�0�u�i�<�(���U���F������e�h�u� ���Gځ�&����W��D^�U���u�u�6�e�j�}����&����V9��T����u�u�u�e�j�}����&����V9��F^�U���u�u�4�1�2�.�W�������lU��h��*���'�&�d�_�w�}�W��������h]��Eߊ�
�
�0�y�w�}�W������F��Q1��F���0�g�"�d�]�}�W���Y���F��Q1��F���0�g�1�y�w�}�W��������h]��Eߊ�
�
�d�n�]�}�W���&����
9��N�����0�!�8��`�l�N���&����Q��1�@���e�u�u�2�9�/�ϳ�	��ƹF�N�����<�!�u�k�d�q�W���Y����W��D�����h�u�y�u�w�}�Wϟ�����d��_N��U���u�u�%�'�w�<�W�ԜY���F��\N��U���6�>�_�u�w�}�W��������E�����u�u�u�1�%�.�G��Y���� 9��1�����&�y�u�u�w�}���D�Ʈ�U9��[����_�u�u�u�w�m�J�������
S��F^�U���u�u�4�1�2�.�W�������l_��h�����d�_�u�u�w�}����Gӄ��lU��W�����u�u�u�u� �l�J�������
S��@����u�u�u�d�j�}����&����WW�N��U���$�u�k�7�1�n�N�������9F���*ي�`�l� �o�4�0����Ӌ��Q��W��E���f�7�3�f�d�h���Y����V��^�����_�u�u�u�w�<�������U��=N��U���u�1�'�&��3���Y��ƹF�N�����&��1�=�j�}�^���YӖ��GF��GN��U���u�u�6�>�j�}�������F�N�����h�u�%�'�#�W�W���Y�ƭ�W��D^��Kʷ�3�f�d�c��9����I���F�N��E��u� �
�
�b�d���s���F�F^��Kʷ�3�f�d�c��m�}���Y���R��R��U��7�3�f�d�a�����
����F�N����h�u� �
��h�N���H���F�N��D��u� �
�
�b�d� ��s���F�S_��Kʷ�3�f�d�c��l�}���Y���BW�	N�����d�c�
�d�l�W�W�������_��h��*���u�:�%�;�9�}�G��L����lV��h]�� ���
�l�d�0�g�}�WϹ�������FךU���u�u�4�4�>�)�W���H���F�N�����&�4�2�u�i�i�}���Y���r��R�����u�k�g�_�w�}�������9F�N��U���u�k�4�
�;�q�W���Y����V��S����&�y�u�u�w�}��������X��B��*��d�0�e�4�3�8���Y���F��R^��Kʷ�3�f�g�f���(���U���F��H��� �
�
�l�f�8�G���U���F������d�h�u� ���N����֓�W��D����u�u�u�0�w�c����J����9��1��D�ߊu�u�u�u�2�}�Iϼ��Փ�
U��R1����_�u�u�u�w�l�J�������_��h��*��_�u�u�u�w�l�J�������_��h��*��n�_�u�u�"��(��H����l3������;�u�e�c�b�l�����Փ�F ��h]�*���_�u�u�0�2�4�W���Y���F�N�����1�=�h�u�e�W�W���Y�ƍ�W��D<�����k�a�_�u�w�}�W�������Z��S�G�ߊu�u�:�!�:�-�_���Y�����S����9�y�u�u�w�}�������R��D�U���u�u�4�1�2�.�W�������lT��1��D���1�0�&�y�w�}�W������F��Q1��G��
�
�
�0�{�}�W���Yӗ��X��B��*��d�0�d�$�{�}�W���YӇ��A��N��U���
�
�l�d�2�l��������9F�N��U���u�k�7�3�d�o�Dށ�&¹��JǻN��U���0�u�k�7�1�n�E��&����D��=N��U���u�d�h�u�"��(��H����l��=N��U���u�d�h�u�"��(��H����l��dךU��� �
�
�c�g�8�G���CӅ��C	��Y��E��`�d�3�e�1�n����J����l��=N��U���0�<�u�4�w�W�W���Y�ƈ�G��S��H���g�_�u�u�w�}����
����T�	N����u�u�u�1�%�.� ������OǻN�����8�%�}�u�w�}�WϽ����R��[�U���u�u�'�&�#�`�W�������F�N�����0�&�u�k�5�;�D��Kù��9��S�����u�u�u�u�4�m�J�������P��h��*���y�u�u�u�w�,�W�������lW��1��E���y�u�u�u�w�<����
�����h]��C���0�e�4�1�2�.�[���Y�����S����f�d�g�
�����Y���F��R_��Kʷ�3�f�d�g���(���U���F�
�H��� �
�
�c�g�8�G���U���F��H��� �
�
�c�g�8�G���P��ƹF��B��*��e�0�d� �m�>��������'��_����3�f�7�3�d�n�B���I�����R��U���u�_�u�u�w�}��������X�BךU���u�u�1�'�$�����D����9F�N��U���'�&��1�?�`�W���Y����\��Z��]���u�u�u�6�<�`�W�������F�N�����!�h�u�%�%�)�}���Y���R��R��U��7�3�f�d�e��(ށ�����@V�N��U���6�e�h�u�"��(��I����l��d��U���u�$�u�k�5�;�D��Kù��9��d��U���u�4�1�0�$�}�Iϼ��Փ�T��R1�����0�&�y�u�w�}�WϽ�H���Q��1�Gڊ�
�
�0�y�w�}�W������F��Q1��D��
�
�
�0�{�}�W���Yӂ��X��B��*��e�0�d�1�{�}�W���Yӗ��X��B��*��e�0�d�$�~�W�W�������l_��h��*���u�:�%�;�9�}�G��L����lV��h]�� ���
�e�
�
�]�}�W�������^��d��U���u��!��3�5�J���K���F�N�����&�4�2�u�i�i�}���Y���r��R�����u�k�g�_�w�}�������9F�N��U���u�k�4�
�;�q�W���Y����V��S����&�y�u�u�w�}��������X��B��*��
�
�
�1�%�.�G�ԜY���F��N��U���
�
�d�
�����Y���F��N��U���
�
�d�
���G�ԜY���F��S�����k�7�3�f�n�m��������@��=N��U���u�0�u�k�5�;�D��I����l��d��U���u�"�d�h�w�(�(܁�Hù��9��BךU���u�u�d�h�w�(�(܁�Hù��9��d��U���u�$�u�k�5�;�D��I����l��dךU��� �
�
�d���(���Y����\��CN��4��d�l�
�
������&����V9��N�����'�6�8�%��}�W���YӢ��R1��C��K��y�u�u�u�w�����
����VF�Z�U���u�u��1�2�.����Y���l�N�����4�u�_�u�w�}�W���Y����C9��\BךU���u�u�0�0�w�c����
��ƹF�N�����&�e�h�u�"��(��&����R��R��Y���u�u�u�6�g�`�W���&����9��1��E�ߊu�u�u�u�g�`�W���&����9��1��Y���u�u�u�4�3�8����Gӄ��lU��^��*ۊ�1�'�&�d�]�}�W���Y����X��B��*��
�
�
�0�{�}�W���Yӑ��[�U��F��e�0�d�"�f�W�W���Y�ƨ�[�U��F��e�0�d�1�{�}�W���Yӗ��X��B��*��
�
�
�d�l�W�W�������U��h��*���u�:�%�;�9�}�G��L����lV��h]�� ���
�e�
�
�]�}�W�������^��d��U���u��!��3�5�J���K���F�N�����&�4�2�u�i�i�}���Y���r��R�����u�k�g�_�w�}�������9F�N��U���u�k�4�
�;�q�W���Y����V��S����&�y�u�u�w�}��������X��B��*��f�0�e�4�3�8���Y���F��R^��Kʷ�3�f�d�f���(���U���F��H��� �
�
�f�d�8�G���U���F������d�h�u� ���D����֓�W��D����u�u�u�0�w�c����J���� 9��1��D�ߊu�u�u�u�2�}�Iϼ��Փ� U��R1����_�u�u�u�w�l�J�������U��h��*��_�u�u�u�w�l�J�������U��h��*��n�_�u�u�"��(��J����l3������;�u�e�c�b�l�����Փ�F ��h]�*���_�u�u�0�2�4�W���Y���F�N�����1�=�h�u�e�W�W���Y�ƍ�W��D<�����k�a�_�u�w�}�W�������Z��S�G�ߊu�u�:�!�:�-�_���Y�����S����9�y�u�u�w�}�������R��D�U���u�u�4�1�2�.�W�������lW��1��D���1�0�&�y�w�}�W������F��Q1��D��
�
�
�0�{�}�W���Yӗ��X��B��*��f�0�d�$�{�}�W���YӇ��A��N��U���
�
�f�f�2�l��������9F�N��U���u�k�7�3�d�l�D܁�&¹��JǻN��U���0�u�k�7�1�n�F��&����D��=N��U���u�d�h�u�"��(��J����l��=N��U���u�d�h�u�"��(��J����l��dךU���!�f�d�m��}�W���	����GF��vX�D���
�
�
�
�"��(��&����F�P�����8�%�}�u�w�}�WϚ�����G�	N�Y���u�u�u��3�8�������R�N��U����1�0�&�>�)�W���K���F��E�����_�u�u�u�w�1�W�������XJǻN��U���0�0�u�k�6����Y���F��S
����h�u�!�f�f�e�(�������l�N��Uʶ�e�h�u�!�d�l�Oׁ���ƹF�N��E��u�!�f�d�o��G�ԜY���F��S�����k�9�
�
�a�e��������9F�N��U���u�k�9�
��k�O���H���F�N��D��u�!�f�d�o����Y���F��N��U���f�d�m�
�f�W�W���Y�ƽ�[�[��*��m�$�|�_�w�}����&����l��h;��U���%�;�;�u�g�k�B���֓�lU��B��*��
�
�_�u�w�8����Y����l�N��Uʑ�!��1�=�j�}�E�ԜY���F��S�����2�u�k�a�]�}�W���Y����V��^
��U��g�_�u�u�8�)����Q���F���U��4�
�9�y�w�}�W�������[�V�����u�u�u�u�6�9����Y����G9��V�*���
�1�'�&�g�W�W���Y�Ư�F���F��a�
�
�
�2�q�W���Y����F���F��a�
�
�
�g�W�W���Y�ƭ�W��D_��Kʹ�
�
�m�c�2�m��������9F�N��U���u�k�9�
��e�A���I����l�N��Uʢ�d�h�u�!�d�l�Cف�&ù��JǻN��U���d�h�u�!�d�l�Cف�&ù��l�N��Uʤ�u�k�9�
��e�A���I����lǻN�����d�a�
�
��}�W���	����GF��vX�D���
�
�
�
�"��(��&����F�P�����8�%�}�u�w�}�WϚ�����G�	N�Y���u�u�u��3�8�������R�N��U����1�0�&�>�)�W���K���F��E�����_�u�u�u�w�1�W�������XJǻN��U���0�0�u�k�6����Y���F��S
����h�u�!�f�f�i�(���&����V��d��U���u�6�e�h�w�)�D��MŹ��9��BךU���u�u�e�h�w�)�D��MŹ��9��d��U���u�4�1�0�$�}�Iϲ�&����P��h_�����&�d�_�u�w�}�W���Y����G9��V�*���
�0�y�u�w�}�Wϩ�H���_��h_�C���d�"�d�_�w�}�W���H���_��h_�C���d�1�y�u�w�}�Wϯ�Y����G9��V�*���
�d�n�_�w�}����L����V9��bN����:�0�!�8��j�F���&ù�� 9��Q1��F���0�e�u�u�0�3�������9F�N��U���4�<�!�u�i�n�[���Y���'��E��'���0�h�u�y�w�}�W���8����@��S��H���|�u�u�%�%�}����s���F�T��H���%�6�>�_�w�}�W�������X��G1���ߊu�u�u�u�3�/���D�Ơ�lU��W�����4�1�0�&�{�}�W���YӅ��[�[��*��`�0�e�6�g�W�W���Y�ƽ�[�[��*��`�0�e�$�{�}�W���YӇ��A��N��U���f�`�l�
������
����F�N����h�u�!�f�b�d�(���&����9F�N��U���u�k�9�
��k�B���I����l�N��Uʱ�u�k�9�
��k�B���I����9F�N��U��h�u�!�f�b�d�(���&���9l�N��*ي�c�`�0�d��g����������Y�Dӳ�e�3�f�7�1�n�D�����ƹF��R �����4�u�_�u�w�}�W�������[F�]����u�u�u�1�%�.�%������JǻN��U���1�'�&��3�5�J���P�����CN�����u�u�u�u�4�6�J���	����l�N��Uʧ�&�!�h�u�'�/��ԜY���F��S�����k�9�
�
�a�h��������@��=N��U���u�0�u�k�;��(��L����l��d��U���u�$�u�k�;��(��L����l��=N��U���u�1�'�&�f�`�W���J����9��1�����&�y�u�u�w�}���D�Ơ�lU��W�����6�d�_�u�w�}�W���Y����G9��X�*���
�0�y�u�w�}�WϺ�Y����G9��X�*���
�d�_�u�w�}�W��D�Ơ�lU��W�����$�|�_�u�w�1�(܁�O�ӓ�lT��T�����;�;�u�e�a�h�Fָ�I����l��h]��Eߊ�
�_�u�u�2�8�������F�N��1����1�=�h�w�o�}���Y���r��R�����u�k�a�_�w�}�W�������@1��C��K��_�u�u�:�#�0����Y���F��[��Kʴ�
�9�y�u�w�}�WϬ�
���F��h��Y���u�u�u�4�3�8����Gӊ�� 9��[��*؊�1�'�&�e�]�}�W���Y����X��C1��@��
�
�
�0�{�}�W���Yӗ��X��C1��@��
�
�
�e�]�}�W���Y����V��S����
�c�`�0�e�<����
��ƹF�N�����k�9�
�
�a�h��������F�N����h�u�!�f�b�d�(���&����9F�N��U��h�u�!�f�b�d�(���&����F�N�����k�9�
�
�a�h��������9F���*ي�m�a� �o�4�0����Ӌ��Q��W��E���f�7�3�f�f�e�}���Y����A��Z��]���u�u�u��#�
����D����l�N��Uʔ�1�0�&�4�0�}�I��s���F�v
�����<�!�u�k�f�W�W�������R�=N��U���u�9�u�k�6����Y���F��R��U��4�
�&�y�w�}�W�������@��
P�� ���
�m�a�4�3�8���Y���F��R^��Kʷ�3�f�d�m��8�[���Y�����
P�� ���
�m�a�$�{�}�W���YӇ��A��N��U���
�
�m�a�6�9����U���F���U��7�3�f�d�o����Y���F��R_��Kʷ�3�f�d�m��8�[���Y�����
P�� ���
�m�a�1�{�}�W���Yӗ��X��B��*��a�$�|�_�w�}��������@��\��*���&�f�
�
�"�1����,�����G�����e�c�`�d�1�m�������� T��h]����
�
� �9�3�-�W�������Z��V�����u�u�u��j�}�[���Y���(��h=��2���k�f�_�u�w�}�W���I����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���:�!����`�W��s���C	����U�ߊu�u�u�u�;�}�IϿ�&����9F�N��U���0�u�k�4��.�[���Y�����N��U���
� �d�g��m�}���Y���W��S����3�
�a�f�'�q�W���Y����C��RN��U���
� �d�g��-����s���F�T��Kʲ�%�3�
�a�d�>�[���Y�����CN��U���
� �d�g��o�L�ԜY�ƪ�9��B��G���f�;�
�g�f�0����	����\��X�����u�e�c�`�f�;�G�������]�� ��F؊�
�4�
�&�]�}�W�������^��d��U���u��u�k�f�W�W���Y�Ƃ�~9��v)��H���y�u�u�u�w�9�߁�0����X�BךU���u�u�<�d� ��?��Y����F�N�����
���u�i�n�^���YӖ��GF��GN��U���u�u�1�;�w�c�������� W��BךU���u�u�<�d�j�}��������9��d��U���u�1� �u�i�:����&����l��dךU���
�
�6�%�d�3�(���
�ד�l3��T�����;�;�u�e�a�h�Fָ�I����C9��Y��G���d�d�u�u�0�3�������9F�N��U���h�u�y�u�w�}�Wϐ�4����t#�	N����u�u�u�<�g�
�3���D����l�N��Uʱ�;�
���w�c�D��Y���F��X��"����h�u�|�w�}����Y����l�N��Uʱ�;�u�k�2�'�;�(��O����9F�N��U���d�h�u�'��(�F��&����F�N�����1�u�k�2�'�;�(��O����\��=N��U���u�:�!�h�w�/�(���H����CT�=d��Uʳ�e�3�8�
�e�.�Dݰ�&¹��fT��N�����0�!�8��`�l�N���&����lU��D1����
�_�u�u�2�8�������F�N��<���k�d�_�u�w�}�W���&����vF�_�U���u�u�1�;���#���G����9F�N��U���d����j�}�E�ԜY���F��B��<���u�k�d�_�w�}�������9F�N��U���e�h�u�8��o����M�ԓ�JǻN��U���<�d�h�u�:��E���&����l��=N��U���u�%�:�0�j�}����K����R��h�����_�u�u�u�w�2���Y����T��B1�A؊�g�n�_�u�w��(���	����@9��Y��*ۊ�g�u�u�:�'�3����I����W��h^�����f�;�
�g�$�l�F���YӁ��V����U�ߊu�u�u�u��`�W��Y���F��b#��!���u�k�d�_�w�}�W����֓�z"��S�F���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���P�����CN�����u�u�u�u�3�3�W�������9��h_�B���y�u�u�u�w�9����GӒ��lQ��Q��A���%�y�u�u�w�}���������hY�����a�b�:�6�3�q�W���Y����\��
P�����`�3�
�a�`�-�^�ԶY����lV��T��Fػ�
�g�&�d�f��C������]����C���d�3�e�3�:��E���J����9��N�����'�6�8�%��}�W���Yӯ��X�d��U���u������J���U���F�
��E�����h�u�e�W�W���Y�ƨ�]W��~*��U��f�y�u�u�w�}����&����{F�_��U���%�'�u�4�w�W�W���Y�ƨ�]V�	N����
� �d�`��m�}���Y���W��S����b�
� �d�b��F�ԜY���F��T��U��!�%�b�
�"�l�B݁�	����l�N��Uʱ� �u�k�!�'�j�(���H����CT�=dװ���u�x�u�=�w�(����Y����VF��G1��*���|�:�u�=�w�)��������VH�d��Uʴ�
��3�8�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W�������l ��R������&�d�3�:�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����Y���F�N��U���u�u�u�%������DӇ��}5��D�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����]	��h����`�<�'�2�f�k�W�������A	��D�X�ߊu�u�'�
�8�8����&����Z9��P1�C܊�&�<�;�%�8�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��M���8�b�|�!�2�}�W���Y���F�N��U���'�
�:�0�#�/�(��&����T9��X��Hʴ�'�;�1�
�2�0�E����ד�V��_����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N�����1�
�0�8�e�h��������F������!�9�g�e�]�}�W���Y���F�R ����u�u�u�u�w�}�������F�N�����<�n�u�u�2�9��������9F�C�ۊ�0�
�f�m�6�.��������@H�d��Uʼ�
�0�
�f�o�<����&����\��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}��������T9��S1�L���!�0�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��Dۊ�&�
�e�|�#�8�W���Y���F�N��U���u�d�'�2�f�j�W������]��[��E�ߊu�u�u�u�w�}�W���������D�����d�l�|�!�2�}�W���Y���F�N��U���d�'�2�d�`�}�JϷ�K����S��h����u�u�u�u�w�}�W���Y����F�N��U���0�1�<�n�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y�ԓ�V��^����2�u�'�6�$�s�Z�ԜY�ƥ�l��h_�E���&�2�
�'�4�g�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��C���8�f�|�u�?�3�}���Y���F�N��U���<�
�0�
�c�m�K���&����T9��]�U���u�u�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y���F�N��G���2�d�e�u�j�<�(���
���� 9��=N��U���u�u�u�u�w�3�W���s���F�N�����<�n�_�u�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������W��V�����'�6�&�{�z�W�W���J����lW��1�����
�'�6�o�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W�������C9��P1����e�|�!�0�w�}�W���Y���F�N��U���'�2�d�d�w�`��������_��UךU���u�u�u�u�w�}����Y�έ�l��D�����
�u�u�%�$�:����&����GU��Q��F���u�=�;�_�w�}�W���Y���F�N��*���
�a�d�i�w��(���&����l�N��U���u�u�u�0�3�4�L���Y���F���U���u�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�4�(���?����\	��D1����m�u�&�<�9�-����
���9F������:�
�:�%�$�/���Aʹ��@��h����%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���J����^9��G�����_�u�u�u�w�}�W���Y���Z*��^1�����:�
�
�0��n�N��Y����Z9��E1�����c�'�2�g�`�f�W���Y���F�N�����u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u�u�u�w�}�;���&����	��h�����f�l�i�u�'�>�����Փ�l�N��U���u�u�u�0�3�4�L���Y���F���U���u�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�4����H����R��P �����&�{�x�_�w�}�(���&����l��^	�����u�u�'�6�$�}������ƹF��R	�����u�u�u�3��-���������������h�r�r�u�?�3�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�W���Y�����R	��F���i�u�
�
�2��D��s���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W�������lW��N�U���6�;�!�9�d�m�}���Y���F�N�����<�n�u�u�w�}�W�������U]�N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ѓ�@��G�����_�u�u�u�w�}�W���Y����]	��h����`�<�d�'�0�o�F���DӇ��l��R1�����d�
�
�
�"�l�G݁�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���f�3�8�f�~�t����s���F�N��U���6�
��������H�ޓ�lV��R	��C���i�u�!�f�f�i�(���&����F�N��U���u�u�6�
���6�������^��h_�����b�e�i�u�#�n�F��&����BV��N��U���u�u�u�u�4��9���8����A��^��*ڊ�0�
�b�`�k�}����H����V9��F_�U���u�u�u�u�w�}����7����a4��E��@ڊ�
�
�0�
�`�m�K����Փ�R��R1����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C�����;�%�:�0�$�}�Z���YӖ��P��F��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y�����Yd��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���������� O������u�u�u�u�w�}�WϽ�&����k'��C��*���
�
�
�0��j�G��Y����lW��1��E���n�u�u�u�w�}�W���YӅ��z(��o/�����
�`�
�
��8�(��L���_��h_�C���d�$�n�u�w�}�W���Y�����~ ��-���!�'�
�`���(���&����Z�[��*��c�0�e�$�l�}�W���Y���F���<�����!�'��h�(���&����Q��R�����
�m�c�0�f�,�L���Y���F�N��U�������#�/�(�������U��S�����d�m�
�d�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���|�!�0�_�w�}�W���Y���F��h��3����:�
�d�2�m����K����[��B��*��f�0�e�$�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�w�}�W���Y���F��[1��*���
�:�%�g���(���&����Z�U��F��e�0�d�$�l�}�W���Y���F�������;� �
�c�o����K����[��d1�� ���;� �
�a�e�;�(��J����9F�N��U���u�u�u�8��o����K����[��Z��G���
�b�b�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�w�}�W���Y���F��[1��*���
�:�%�g���(���&����Z�U��F��g�
�
�
�g�W�W���Y���F�N��*����'��:��j��������R��S�� ���
�c�e�0�f�,�L���Y���F�N��U���
�8�d�
��8�(��H���@��C��D���3�
�l�l�'�f�W���Y���F�N�����8�g�
�
�2��A��E�ƿ�_9��G\�����
�e�f�%�l�}�W���Y���F���*���g�
�
�0��k�D��Y����G��1�����e�d�%�n�w�}�W���Y���F��R����
�
�0�
�a�d�K�������CU��^1��*��b�%�n�u�w�}�W���Y�����hY�����g�`�u�h�#�-�@ہ�����9��d��U���u�u�u�u�w�)���&����P��R�����m�
� �d�a��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��B���8�g�|�|�#�8�}���Y���F�N�����!��'��8��B���I����lT��N�U���
�
�l�d�2�m���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Fڊ�&�
�l�|�w�5����Y���F�N��U�������#�h�(���&����Z�Q=��0���� �
�c�1��@���	��ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z���
������T��[���_�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�n�t�W������F�N��U���u��-� �.�(�(�������R��S����� �d�g�
�e�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l�� 1����|�|�!�0�]�}�W���Y���F�^"�����'��:�
�a�/���N�����[�����:�%�d�
�"�l�Cց�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�)��ԜY���F�N��Uʼ�d�'�2�g�o�}�JϷ�H����R��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�n�(���&���F��R ךU���u�u�u�u�w�}�(܁�����U�
N��F���
�d�b�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�w�}�W���Y���F��hZ�����b�f�i�u�����MŹ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��E������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���|�u�=�;�w�}�W���Y���F��R	��A��i�u�'�
�"�l�E܁�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�a�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��]��\���=�;�u�u�w�}�W���Y����V��X�I���'�
� �d�d��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Fي�&�
�g�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&���� U�G�����u�u�u�u�w�}�W�������Q��S�����d�m�
�e�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���4�1�}�%�4�3����H�����C��؊� �d�a�
�e�t�W������F�N��U���u�8�
�d�%�:�E��Q���F��G1�*���d�`�
�d�g�f�W�������9��P1�M���|�i�u�8��l����L�ӓ�N��d��Uʡ�%�f�
�0��i�F��Y����^��1��*���`�%�}�|�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��Q��F���4�1�}�%�4�3����H�����C��ۊ� �g�g�
�e�t�W������F�N��U���u�8�
�a�%�:�E��Q���F��G1�*���g�f�
�d�g�f�W�������9��P1�C���|�i�u�8��i����H�Փ�N��d��Uʡ�%�f�
�0��j�O��Y����^��1��*��f�%�}�|�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��Q��F���4�1�}�%�4�3����H�����C�����
�d�e�%�~�t����s���F�N��U���!�%�f�
�2��@��I�����h]�����d�g�%�}�~�W�W�������l��h\�M��u�h�!�%�d����L����W�=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�g�1�0�F�������K��X ��*���d�b�
�g�j�<�(���
����9��G�����u�u�u�u�w�}�W�������V��W�E���h�!�%�3��i�N���Q����F�C�����g�l�}�|�k�}��������
9��_����u�8�
�0��n�G��Y����^��B1�Mӊ�d�g�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=N��U���
�
�`�
�3�/����K����F��@ ��U���i�u�e�w�]�}�W���&����_��S
�����g�c�}�u�8�3���Y���V�=N��U���f�d�m�
�3�/����K����F��@ ��U���i�u�e�w�]�}�W���&����R��S
�����g�b�}�|�k�}�G��Y����^��R	��F��c�u�:�;�8�n�W��[����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ƹ�C9��h��*��d�c�u�:�9�2�D���D����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G���s���G��Z�����b�m�c�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��[���F��G1�*���
�b�m�c�w�2����K���D��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I���9l�N�U���u�0�!�&�6�8�_���7����^O��QN��ʦ�4�0�8�6�>�8�W��Y����C9��h��*���<�;�%�:�w�}����
����C9��V��U����
�&�y�6���������V��h�����4�
� �g�g�-�[ϻ�����WS��B1�B݊�g�u�-�!�8�9�(���H����CT�R�����f�3�
�`�c�-�[ϻ�����WT��B1�Aي�g�u�-�!�8�9�(���K����CT�R�����
� �g�a��o�}���Y����]l�N��Uʶ�&�u�%���.�W���Y���F�N�����4�
��&�f�;���D��ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u���������T�����2�6�e�|�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��D�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����]��QUךU���u�u�u�u�?�3����-����l ��h_��K�ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��^�����3�
�a�b�'�}�W�������l
��h^��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�C�������F�N��U���u�u�0�&�1�u�_�������l
��^��U���%�6�|�4�3�u��������U��Y�����u�%�6�;�#�1�F��P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��[��U���u�u�u�u�w�}�W�������l ��R������&�g�3�:�l�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��F���8�g�h�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�d�;���s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���a�3�8�f�j�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!��.�(��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�C�������F�N��U���u�u�0�1�>�f�W���Y���F��_������&�`�3�:�i�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���L����lR��N��U���u�u�u�u�2�9���Y���F�N�����4�
��&�a�;���D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����l ��h[�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�@������FǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3����	����@��A_��U���-�!�:�1��(�F��&���O��_��U���u�u�u�u�w�}�W�������l ��R������&�l�3�:�e�}���Y���F�N�����3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)����I����K��X ��*���d�l�
�g�~�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��B���8�c�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����9��Z1�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���m�3�8�b�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���e�3�8�l�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:�����3�8�l�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�d�1�0�F��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�F߁�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�d�1�0�F���G���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	���&����W��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����W��D��E�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���K����lW��
P��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]9��D��E���4�
�0�1�1��N߁�K����C9��Y�����e�|�4�1��-��������lV������1�
� �d�e��E���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�d�n�w�}�W���Y���F��[��U���4�
�:�&��2����Y�ƭ�l����U���;�'�&�!�g�/��������F9��1��U���%�6�;�!�;�l�G���ӈ��N��h�����#�
�u�u�/�)����&����T��G\��\���!�0�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	���&����T�	NךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�d�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��1����u�k�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�c�W�W���Y���F�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�c�;���B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�`�3�8�f�}�I�ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$����ӓ�@��UךU���u�u�u�u�w�}�������F�N��Uʢ�0�u�%���)�A�������X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�
���F�N��U���u�u�u�4������E�ƭ�l5��D�*���
�`�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����Q��D��C��u�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	�������!�9�d�e�j�8�����ԓ�F9��]��G���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���J����lU��=N��U���u�u�u�u�w�1����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[��E��0�<�6�;�e�;�(��J����O��_��U���u�u�u�u�w�}�W�������l ��R������&�d�
�$��@�ԜY���F�N��Uʰ�&�_�u�u�w�}�W���Y���F��h �����i�u�%���)�@�������9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�m�1�0�F���G���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	���&����^��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����^��D��B�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���@����lW��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�m�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��^�����l�h�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���7����^F���&���!�d�3�8�e�f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�e�����@���F�N��U���u�0�1�<�l�}�W���Y�����YN��*���&�g�
�&��m�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�E�������9F�N��U���u�u�u�9�2�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��^�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�E݁�
����[�=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����U��D��G�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��G���8�g�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GT��Q��G���k�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�f�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�f�1�0�E��Y���F�N��U���;�u�3�_�w�}�W���Y�ƻ�V��G1��*���a�3�8�g�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�e�����M���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���M����lT��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�h����K���l�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��[�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��[�����a�_�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�"�2�}����&����l ��h\�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��B���8�g�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�g�
�&��h�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��G݊�&�
�c�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�m�1�0�E��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�E؁�
����l�N��U���u�u�u�0�3�4�L���Y���F���ʴ�
��&�g��.�(��D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���@����lT��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GT��Q��G��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���Kʹ��^9��S����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�4�
��;���Y����g9��^�����l�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���l�3�8�g�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӈ��`2��C]�����g�u�k�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�f�
�&��m�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�m����K��ƹF�N��U���u�u�;�u�1�W�W���Y���F��R �����
�!�d�3�:�n�W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�D݁�
����l�N��U���u�u�u�0�$�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����l ��h]����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��D��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��F؊�&�
�d�_�w�}�W���Y���F��SN��N���u�u�u�u�w�*����	����@��h��*��h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���a�3�8�f�l�}�W���Y���F������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�f��.�(��s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���f�
�&�
�d�`�W���Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�h����J��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���Jǹ��^9��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���;�4�
��$�n�(���&���FǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3����	����@��A_��U���-�!�:�1��(�E��&���O��_��U���u�u�u�u�w�}�W�������l ��R������&�f�
�$��A�ԜY���F�N��Uʰ�&�3�}�}�'�>��������lW������4�1�}�%�4�3����H�����C��ۊ� �g�g�
�e�t�W������F�N��U���u�u�u�%������DӇ��`2��C]�����f�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���f�
�&�
�c�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�`�h�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�`�3�:�n�L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�n�(���&����F�N��U���u�u�0�1�>�f�W���Y���F��_������&�f�
�$��A��Y���F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��-��������lV������1�3�
�d�g�-�^���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ۊ�&�
�n�u�w�}�W���Y�����^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�#��}�W�������l ��_�*��|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���J˹��^9��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$����ޓ�@�� N��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�%������DӇ��`2��C]�����f�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���f�
�&�
�`�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƣ�[��S�U���u�u�u�u�w�}�WϿ�&����@�
N��-���������/���!����k>��o6��-���w�_�u�u�w�}��������F�R �����0�&�_�u�w�p�W�������R��P �����&�{�x�_�w�}��������@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}����UӇ��@��T��*���&�f�
�&��k�W�������l ��_�*��_�u�u�0�>�W�W���Y�ƥ�N�Y��]���6�;�!�9�0�>�F������R��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��X�����;�!�}�%�4�3����H�����C�����
�d�e�%�~�t�^Ϫ���ƹF�N��U���%�1�;�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��X ��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���0�4�&�2�w�/����W���F�V�����4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�N�����;�u�u�u�w�4�W�������C9��Y�����6�d�h�4��)����Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�]�}�W���Y���R��S��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������R��V�����'�6�&�{�z�W�W���	����W��D�����:�u�u�'�4�.�_�������C9��P1������&�f�
�$��A�������]��B1�Aڊ�g�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��B���8�f�|�4�3�3����	����@��A_��U���-�!�:�1�1��F���	���F��R ��U���u�u�u�u�6�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�0�1�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�%�'�!�%��W������w#��e<�����a�
�
�
�2��A��s���R��R����i�u�9����%�������9��1����e�n�u�u�6��������F��h'��0����0�8�d�g�8�G�������]ǻN�����!�'�
�u�j�>�(���<����G��h_�*���
�0�
�b�g�W�W���	����F��N�U�������#�/�(��&����A��Y�N���u�4�
�0�"�3�B��Y����}"��v<�����d�g�0�d�%�:�E��B�����E�����u�h�6�
���6�������R��h^�����b�e�_�u�w�-��������[��[1��1����!�'�
�b��(ށ�����S��N�����0� �;�m�k�}����M����F�V�����;�l�i�u���3���+����^9��h��*��`�_�u�u�z�}��������lW�������%�:�0�&�w�p�W�������T9��S1�M���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�m�i�w�<�(���
����9��
N��*���3�8�g�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��]����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��l�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�d�d�}�J���	����@��A_��U���%��
�&��e��������O��N�����%�:�0�&�]�W�W���TӇ��@��U
��D��4�&�2�u�%�>���T���F��h��*���
�c�
�&�>�3����Y�Ƽ�\��DF��*���3�8�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��k�W��Q����\��h��*���u�%��
�$�u�AϺ�����P�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����m�4�&�2�w�/����W���F�V�����1�
�b�
�$�4��������C��R������3�8�_�w�}����s���F�N��U���4�
�<�
�3��@���D�έ�l��D��ۊ�u�u�%���.�_������\F��G�U���0�1�%�:�2�.�}�ԜY�����D�����d�l�4�&�0�}����
���l�N��*���
�1�
�m��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��Y���R��X ��*���
�u�u�%������Kӂ��]��\��N���u�0�1�%�8�8��Զs���K��G1�����1�d�l�u�$�4�Ϯ�����F�=N��U���&�2�7�1�f�d�(�������A	��N�����&�4�
�0�w�3�����֓�V��E��*���g�e�%�|�w�}�������F�N��U���u�%�&�2�5�9�F��Y�����T�����2�6�d�h�6������Ƣ�GN��Y1�����e�'�4�
�2�9����@ù��[��G1�����9�d�e�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@�ƭ�@�������{�x�_�u�w�-��������_��V�����'�6�o�%�8�8�ǿ�&����P��h=����
�&�
�d�w�%��������lW��1��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�l�u�j�u��������_	��T1�Hʴ�
�<�
�&�&��(���K����lW����U´�
�:�&�
�!��W�������]��Q��@���%�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�l�G���
������T��[���_�u�u�%�$�:����H����R��P �����o�%�:�0�$�<�(���&����l5��D�*���
�a�u�-�#�2�ށ�����9��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����e�u�h�}�6�����&����P9��
N��*���
�&�$���)�B��������� ��]´�
�:�&�
�!��W�������]��Q��D���%�|�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��N���
������T��[���_�u�u�%�$�:����H�ѓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��Y��H���%�6�;�!�;�l�F������l ��]����!�u�f�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z�F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�3����	����A������!�9�2�6�g�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����g�i�u�4��2����¹��F��h-�����d�1�"�!�w�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����a�i�u�4��2����¹��F��h-�����c�1�"�!�w�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����l�i�u�4��2����¹��F��h-�����d�u�:�;�8�l�^��Y����]��E����_�u�u�x�w�-��������W��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��Z�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����f�d�i�u�6�����&����F�V��&���8�d�u�:�9�2�F���B����������n�_�u�u�z�}��������lU�������%�:�0�&�w�p�W�������T9��S1�F���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�f�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��[�����;�%�:�0�$�}�Z���YӇ��@��U
��F���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�f�`�k�}��������_��N������3�8�d�w�2����H���9F���U���6�&�n�_�w�}�Z���	����l��h]�U���<�;�%�:�2�.�W��Y����C9��P1����b�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�f�`�a�Wǿ�&����G9��1�Hʴ�
��3�8�f�}��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��E���&�<�;�%�8�8����T�����D�����a�m�4�&�0�����CӖ��P����6���&�|�u�u�5�:����Y���F�N��U���&�2�7�1�c�e�K�������]��[��D��4�
��3�:�l�W������O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�a�e�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�i�G��Yۇ��P	��C1��D��h�4�
��1�0�F�������W��UךU���;�u�'�6�$�f�}���Y���R��^	�����f�u�&�<�9�-����
���9F������7�1�a�d�6�.���������T��]����
�&�|�w�}�������F�N��U���u�%�&�2�5�9�C��E����C9��Y�����d�h�4�
��;���Y����G	�G����u�;�u�'�4�.�L�ԶY���F��h��*���
�a�u�&�>�3�������KǻN�����2�7�1�a�f�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���H�����T�����d�d�h�4������K�ƨ�D��\�\�ߊu�u�;�u�%�>���s���K�V�����1�
�`�u�$�4�Ϯ�����F�=N��U���&�2�7�1�c�d��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����M���F��G1�����9�d�d�h�6��$�������W	��C��A���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�c�w�.����	����@�CךU���%�&�2�7�3�i�N���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(������F��@ ��U���|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�o�}����Ӗ��P��N����u�%�&�2�5�9�C�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������U�
N�����;�!�9�d�f�`����*����T��S�����m�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��d�W�������A	��D�X�ߊu�u�%�&�0�?���O����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lR��R��]���6�;�!�9�f�l�JϿ�&����@�N�����u�l�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��F���
������T��[���_�u�u�%�$�:����L�֓�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��^��H���%�6�;�!�;�l�F������l ��]����!�u�e�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(������]F��X�����x�u�u�4��4�(���&�Г�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U´�
��3�8�g�9� ���Y�����T�����d�d�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�h�GϿ�
����C��R��U���u�u�4�
�>�����Où��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��Z�����:�f�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�B������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��V�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�f�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���AӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�M��u�4�
�:�$��ށ�Y�ƭ�l%��Q��Gʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@Ӈ��Z��G�����u�x�u�u�6���������
9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�4�
�:�$��ށ�Y�ƭ�l%��Q��@ʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���NӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�B��u�4�
�:�$��ށ�Y�ƭ�l%��Q��Bʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@Ӈ��Z��G�����u�x�u�u�6���������
9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�4�
�:�$��ށ�Y�ƭ�l%��Q��D���:�;�:�d�~�f�W�������A	��D����u�x�u�%�$�:����A����@��YN�����&�u�x�u�w�<�(���&����Q��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��M��i�u�4�
�8�.�(���&���R��d1����u�:�;�:�f�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����m�i�u�4��2����¹��F��h-�����f�u�:�;�8�n�^��Y����]��E����_�u�u�x�w�-��������^��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��V�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����m�m�i�u�6�����&����F�V��&���8�f�u�:�9�2�D���B����������n�_�u�u�z�}��������l^�������%�:�0�&�w�p�W�������T9��S1�M���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�m�m�i�w�<�(���
����9��
N��*���3�8�f�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��[�����;�%�:�0�$�}�Z���YӇ��@��U
��L���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�l�`�k�}��������_��N������3�8�f�3�*����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��[�����;�%�:�0�$�}�Z���YӇ��@��U
��L���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�l�`�k�}��������_��N������3�8�a�3�*����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��Y�����;�%�:�0�$�}�Z���YӇ��@��U
��L���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�l�b�k�}��������_��N������3�8�m�3�*����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��^�����;�%�:�0�$�}�Z���YӇ��@��U
��L���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�l�e�k�}��������_��N������3�8�l�3�*����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��[�����;�%�:�0�$�}�Z���YӇ��@��U
��L���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�l�`�k�}��������_��N������3�8�g�w�2����K���9F���U���6�&�n�_�w�}�Z���	����l��F1��*���e�3�8�l�6�.��������@H�d��Uʴ�
�<�
�&�&��(���I����l_��D�����:�u�u�'�4�.�_���
����W��^��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��L��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�e�3�:�d�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�l�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�d�3�8�f�}����Ӗ��P��N����u�%�&�2�4�8�(���
����U��^�����;�%�:�u�w�/����Q����Z��S
��@���u�u�7�2�9�}�W���Yӏ����D�����m�l�u�=�9�W�W���Y���F��h��*���$��
�!�f�;���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���H����lW��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!�e�;���Y����T��E�����x�_�u�u�'�.��������l��1����
�&�<�;�'�2�W�������@N��h��*���
�d�|�u�w�?����Y���F��QN�����2�7�1�f�n�}����s���F�N�����<�
�&�$����������F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����T��D��D��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$����������F��D��U���6�&�{�x�]�}�W���
����@��d:�����3�8�d�
�$�4��������C��R�����<�
�1�
�c�t�W�������9F�N��U���}�%�&�2�5�9�D��Y����l�N��U���u�4�
�<��.����&����l ��h_�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(���&����l5��D�*���
�g�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��.����&����l ��h_����2�u�'�6�$�s�Z�ԜY�ƭ�l��h�����
�!�a�3�:�l�(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��Z�����f�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���d�
�&�
�d�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9��[�����a�4�&�2�w�/����W���F�V�����&�$��
�#�h����Hǹ��@��h����%�:�0�&�6���������OǻN�����_�u�u�u�w�;�_���
����W��[�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�a�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�d��.�(��E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�`�6�.��������@H�d��Uʴ�
�<�
�&�&��(���O����lW��V�����'�6�o�%�8�8�ǿ�&����Q��Y����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�d�
�$��B��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�Fف�
����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�d�
�$��AϿ�
����C��R��U���u�u�4�
�>�����*����Q��D��C���&�2�
�'�4�g��������C9��P1����b�_�u�u�2�4�}���Y���Z �V�����1�
�b�|�#�8�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
����U��X��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�l�(���&����@��YN�����&�u�x�u�w�<�(���&����l5��D�*���
�b�4�&�0�����CӖ��P�������7�1�a�m�]�}�W������F�N��U´�
�<�
�1��m�^Ϫ���ƹF�N��U���%�&�2�6�2��#���H˹��^9��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���Hʹ��^9�������%�:�0�&�w�p�W�������T9��R��!���d�
�&�
�o�<����&����\��E�����%�&�2�7�3�l�D���Y����V��=N��U���u�3�}�%�$�:����H������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���l�3�8�d�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��h��*���&�<�;�%�8�8����T�����D�����
��&�d�1�0�G���
����C��T�����&�}�%�&�0�?���P�����^ ךU���u�u�3�}�'�.����������YNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:��ۊ�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����9��Z1�U���<�;�%�:�2�.�W��Y����C9��P1������&�g�
�$��N���
����C��T�����&�}�%�&�0�?���I���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��C\�����d�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�e�3�8�f�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C\�����g�u�&�<�9�-����
���9F������6�0�
��$�o�(���&�֓�@��Y1�����u�'�6�&��-�������� W�N�����;�u�u�u�w�4�Wǿ�&����Q��]�U���;�_�u�u�w�}�W���	����l��F1��*���d�3�8�g�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!�f�;���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���g�3�8�g�w�.����	����@�CךU���%�&�2�6�2��#���K����^9��h�����%�:�u�u�%�>����	����l��hZ�\���u�7�2�;�w�}�W�������C9��P1����d�u�=�;�]�}�W���Y���R��^	������
�!�g�1�0�E���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$����������F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�f�1�0�E���
������T��[���_�u�u�%�$�:����&����GT��Q��G؊�&�<�;�%�8�}�W�������R��^	�����`�|�u�u�5�:����Y����������7�1�d�m�w�5��ԜY���F�N��*���
�&�$���)�D�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����l ��h\�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�C�������R��P �����&�{�x�_�w�}��������B9��h��A���8�g�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�b�~�}�Wϼ���ƹF�N�����%�&�2�7�3�l�O������F�N��U���4�
�<�
�$�,�$����ғ�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��Z�����f�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����ӓ�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�`�3�8�e���������PF��G�����4�
�<�
�3��B���Y����V��=N��U���u�3�}�%�$�:����M���G��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�a�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*���4�&�2�u�%�>���T���F��h��*���$��
�!�a�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lR��N�����u�u�u�u�w�}��������V��c1��G܊�&�
�`�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�g�
�$��B��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��G݊�&�
�c�4�$�:�W�������K��N�����<�
�&�$����������9��D��*���6�o�%�:�2�.��������W9�� GךU���0�<�_�u�w�}�W���Q����Z��S
��C���!�0�u�u�w�}�W���YӇ��@��T��*���&�g�
�&��k�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�o�(���&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�g�
�&��j�����Ƽ�\��D@��X���u�4�
�<��.����&����l ��h\�����2�
�'�6�m�-����
ۇ��@��U
��L���_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�l�|�!�2�}�W���Y���F��G1�����0�
��&�e�����N���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���K˹��^9��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�e�����AӇ��Z��G�����u�x�u�u�6�����
����g9��W�����m�4�&�2��/���	����@��G1�����1�a�f�_�w�}����s���F�^�����<�
�1�
�o�t����Y���F�N��U���&�2�6�0��	���&����^�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����GT��Q��G���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��G���8�d�4�&�0�����CӖ��P�������7�1�g�g�]�}�W������F�N��U´�
�<�
�1��e�^Ϫ���ƹF�N��U���%�&�2�6�2��#���K����lW�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����GT��D��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�D߁�
������^	�����0�&�u�x�w�}��������V��c1��Fڊ�&�
�l�4�$�:�(�������A	��D�����2�7�1�a�a�W�W�������F�N�����4�
�<�
�3��N�������9F�N��U���u�%�&�2�4�8�(���
����U��W��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C]�����g�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��^�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�f�
�&��m��������\������}�%�&�2�5�9�B��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���d�3�8�f�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�d�����H����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�f�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�g�1�0�D���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:�����3�8�f�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	���&���� T��D�����:�u�u�'�4�.�_���
����W��W��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��D��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�f�3�:�n�W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�D�������[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��h�����
�!�a�3�:�n�W�������A	��D�X�ߊu�u�%�&�0�>����-����9��Z1�*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�d�b�u�?�3�}���Y���F�V�����&�$��
�#�i����J�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$����ғ�@��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�h����J�ƭ�@�������{�x�_�u�w�-��������`2��C]�����f�
�&�<�9�-����Y����V��V�����1�
�c�|�w�}�������F���]���&�2�7�1�b�m�W������F�N��Uʴ�
�<�
�&�&��(���L����lU��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���O����lU��V�����'�6�&�{�z�W�W���	����l��F1��*���c�3�8�f��.����	����	F��X��´�
�<�
�1��e�^���Yӄ��ZǻN��U���3�}�%�&�0�?���A�Ƹ�V�N��U���u�u�4�
�>�����*���� P��D��@��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��F܊�&�
�`�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�>�����*���� Q��D��Cʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�b�1�0�Dف�
����l��TN����0�&�4�
�>�����A��ƹF��R	�����u�u�u�3��-��������W�C��U���u�u�u�u�w�<�(���&����l5��D�*���
�c�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�f�
�&��k�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�*���
�b�4�&�0�}����
���l�N��*���
�&�$���)�O�������R��P �����o�%�:�0�$�<�(���&����_��=N��U���<�_�u�u�w�}����	����l��hV�\ʡ�0�u�u�u�w�}�W�������T9��R��!���f�
�&�
�`�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�d�����N���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���f�3�8�g�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&����9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��G���!�0�u�u�w�}�W���YӇ��@��T��*���&�f�3�8�e�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�d�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=�����3�8�f�4�$�:�W�������K��N�����<�
�&�$���ہ�
����R��P �����o�%�:�0�$�<�(���&����
W��=N��U���<�_�u�u�w�}����	����l��hW�\ʡ�0�u�u�u�w�}�W�������T9��R��!���a�3�8�f�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�a�1�0�D��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��@���8�a�4�&�0�}����
���l�N��*���
�&�$���)�(���&ǹ��@��h����%�:�0�&�6���������OǻN�����_�u�u�u�w�;�_���
����W��[�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�a�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�`�3�:�i�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�����`�4�&�2�w�/����W���F�V�����&�$��
�#�����&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������l^��N�����u�u�u�u�w�}��������V��c1��C���8�`�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�c�3�8�b�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9�� 1����4�&�2�u�%�>���T���F��h��*���$��
�!��.�(ف�
����l��TN����0�&�4�
�>�����I��ƹF��R	�����u�u�u�3��-��������R�C��U���u�u�u�u�w�<�(���&����l5��D�����c�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���b�3�8�c�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��Q��Bʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�
�$��(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��1����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�b�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�>�����*����
9��Z1����2�u�'�6�$�s�Z�ԜY�ƭ�l��h�����
�!�
�&����������PF��G�����4�
�<�
�3��C���Y����V��=N��U���u�3�}�%�$�:����@���G��d��U���u�u�u�4��4�(�������@��Q��M��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��L���8�m�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʴ�'�;�1�
�2�0�E����ד�F9��\��G��u�!�
�:�>�����ۓ��Z��SF�����1�
�0�8�e�h��������O������1�4�
�:�$��݁�P��ƹF��B��*��f�0�e�4�3�8����DӒ��lU��E��G��}�u�u�u�8�3���B���F���*ي�f�f�0�e�6�9����Y����T��E�����x�_�u�u�"��(��J����l��E��D���&�2�
�'�4�g��������C9��P1������&�d�
�$��E���	����l��F1��*���a�3�8�d�{�<�(���&����l5��D�*���
�a�u�%�$�:����&����GW��Q��D���u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�u�=�9�W�W���Y���F��Q1��D��
�
�
�1�%�.�F��Y����\��h��A��g�x�d�1� �)�W���s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�`�3�:�l�^������F�N��U���7�3�f�d�d��(߁�����@W�
N��*���&�
�#�a�e�o�Z������\F��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���������� O�C��U���u�u�u�u�w�?����H����V9��V
�����u�h�4�
�8�.�(���M���K�
�����e�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y����F ��h_�F���e�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����RNךU���u�u�u�u�"��(��J����l��E��D��u��w�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y���� 9��]��*ڊ�0�u�&�<�9�-����
���9F���*ي�f�f�0�e�4�m��������\������}�%�6�y�6�����
����g9��Z�����f�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��A���8�g�|�|�#�8�W���Y���F���*ي�f�f�0�e�4�m�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���*ي�f�f�0�e�4�m�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����H����V9��T����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��]�*���
�0�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��\����<�
�&�$���������� J��G1�����0�
��&�f�����M�ƭ�l��h�����
�!�c�3�:�l�^���Yӄ��ZǻN��U���3�}�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�d�;���P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��Z�����f�|�:�u��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��C���8�d�|�|�w�5��ԜY���F�N�����d�f�
�
��8�W������]��[����_�u�u�u�w�1��ԜY���F�N�����d�f�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�"��(��J����l��S�� ���
�e�
�
��m�}���Y���Q��1�Fي�
�
�0�u�$�4�Ϯ�����F�=N��U���
�
�f�f�2�m� �������]9��X��U���6�&�}�%�4�q��������V��c1��Dي�&�
�g�u�'�.��������l��1����y�4�
�<��.����&����l ��h_�U���&�2�6�0��	���&����S�N�����;�u�u�u�w�4�W���Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��\��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�a�3�:�l�^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����S��D��A���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��P����[��=N��U���u�u�u� ���D����֓�VW�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u� ���D����֓�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���Yӄ��lU��]�����4�1�0�&�w�`����J¹��T9��_��U���u�:�;�:�g�f�}���Y����F ��h_�F���d�4�1�0�$�}����Ӗ��P��N����u� �
�
�d�n��������@��V�����'�6�o�%�8�8�ǿ�&����P��h=����
�&�
�g�w�-��������`2��C_�����d�y�4�
�>�����*����S��D��A���%�&�2�6�2��#���HŹ��^9��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���� 9��]��*ۊ�1�'�&�d�k�}��������EP��F�X��1�"�!�u�~�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N�����d�f�
�
��9����H���R��X ��*���a�g�g�x�f�9� ���Y����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!�c�;���P�Ƹ�V�N��U���u�u�7�3�d�l�D܁�&¹��W��D_��Hʴ�
�:�&�
�!�i�F��T����\��XN�N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����Փ�@��G�����u�u�u�u�w�}�Wϼ��Փ� U��R1�����0�&�u�h�6�����&����lV�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�d�n��������@��S��-���_�u�u�u�w�3�W���Y����������n�_�u�u�z�}����&����l��h��U���<�;�%�:�2�.�W��Y����F ��h_�F���d�6�e�4�$�:�(�������A	��D�����y�4�
�<��.����&����l ��h_����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��Q��D���|�!�0�u�w�}�W���Y����F ��h_�F���d�6�e�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����F ��h_�F���d�6�e�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�7�3�d�l�D܁�&¹��F��D��U���6�&�{�x�]�}�W���&���� U��h_��ۊ�&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�F܁�
����F��h��*���$��
�!�c�;���UӇ��@��T��*���&�d�
�&��i�W���
����@��d:�����3�8�d�|�w�}�������F���]���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�f�3�8�f�t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��C������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�u�=�;�]�}�W���Y���Q��1�Fي�
�
�0�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���Q��1�Fي�
�
�0�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u� �
�
�d�n���������h]��Eߊ�
�
�e�_�w�}�Z�������U��h��*���u�&�<�;�'�2����Y��ƹF��B��*��f�0�d�"�f�<����&����\��E�����%�6�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
����U��]����<�
�&�$����������J��G1�����0�
��&�f�����L���F��P��U���u�u�<�u��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�F܁�
����O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���L����lW��N��U���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�b�t�^Ϫ���ƹF�N��U��� �
�
�f�d�8�F���H���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U��� �
�
�f�d�8�F���H���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����J����
9��S����� �a�m�%�w�`��������_��h^��U���u�:�;�:�g�f�W�������lW��1�����&�u�h�!�'�n�(���H����CW�C��U���;�:�e�n�]�}�W������lW��1�����&�u�&�<�9�-����
���9F���*ي�`�l�4�1�2�.�(�������A	��N�����&�7�3�f�f�k�(�������lT�� B�����2�6�0�
��.�E������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�f�u�:��N���&����l��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����U�� G�����u�u�u�u�w�}�Wϼ��Փ�P��V
�����u�h�!�%�e����Hʹ��T�_�����:�e�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y����F ��h_�L���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��G���8�d�|�!�2�}�W���Y���F��B��*���l�4�1�0�$�}�Jϼ��Փ�P��V
��*���
�f�b�_�w�}�W������F�N��U���7�3�f�d�a�����
���F��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�n�F��&����R��P �����&�{�x�_�w�}����&����l��h�����%�:�u�u�%�>����	������D�����
��&�d��.�(��s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�j����H�����YNךU���u�u�u�u�"��(��@����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u� �
��h�N���I���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������lW��1��Dʴ�&�2�u�'�4�.�Y��s���Q��1�Cӊ�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K����lW�V�����&�$��
�#�����UӇ��@��T��*���&�a�3�8�d�W�W�������F�N�����}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�^ϱ�Y�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��hY��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^������F�N��U���7�3�f�d�a�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����f�d�c�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�(�(܁�L�ߓ�F��D��U���6�&�{�x�]�}�W���&����_��1�����
�'�6�o�'�2��������lW��h^�����d�0�d�w�?�D��L����F��h��*���$��
�!��.�(������T9��R��!���m�3�8�b�w�-��������`2��CZ�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��Q1��D��
�d�i�u�5�n�F��&����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�7�3�f�f�k�(��E�ƥ�l5��1��D�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ԓ�@��G�����_�u�u�u�w�}�W���&����_��N�U����
�
�
�l�}�W���YӃ��VFǻN��U���u�u� �
��h�N���Y���k>��o6��-���������/���!����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���7�3�f�d�a�����
������T��[���_�u�u� ���B����ד�@��Y1�����u�'�6�&��-�������T9��R��!���g�3�8�d�w�%����ƹ��lW�� 1��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�c�;���s���Q��Yd��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�e����N����AF�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����|�4�1�;�#�u��������U��Y�����u�%�6�;�#�1�F��P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�|�!�0�w�}�W���Y�����h]��@���"�d�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���Yӄ��lU��X����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N�����d�g�
�
��9����I���G��_�����a�d�g�x�f�9� ���Y����9F�C����f�d�g�
������
����@��YN�����&�u�x�u�w�?����H����V9��V
�����
�&�<�;�'�2�W�������@N��h��*���$��
�!��.�(������T9��R��!���d�
�&�
�g�}��������B9��h��*���
�y�4�
�>�����*����V��D��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���Q��1�Gڊ�
�
�1�'�$�l�K���	����@��AX��F��x�d�1�"�#�}�^�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�t����Y���F�N��U���
�
�c�e�2�m��������[��G1�����9�c�
�}�w�}�W������]ǻN��U���9�<�u�}�'�>��������lW������6�0�
��$�d����A����[��=N��U���u�u�u� ���A����֓�W��D�I���%�6�;�!�;�k�(���Y����W	��C��\�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ѓ�@��G�����_�u�u�u�w�}�W���&����V��h^�����&�d�i�u�'�>��������N��N����!�u�|�_�w�}�W������F�N��U���7�3�f�d�e��(߁�����@W�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����H����V9��T����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��X�*���
�0�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��W��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� V��D��L���u�=�;�_�w�}�W���Y�Ʈ�U9��X�*���
�0�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ʈ�U9��X�*���
�0�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u� �
��k�G���I������^	�����0�&�u�x�w�}����J����9��1��D���&�2�
�'�4�g��������C9��N��*���
�&�$���)�(���&����C9��P1������&�d�
�$��G���	����l��F1��*���
�&�
�y�6�����
����g9��^�����|�u�u�7�0�3�W���Y����UF�F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�F�������F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��L���8�m�|�:�w�u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�F߁�
����O�C��U���u�u�u�u�w�?����H����V9��T�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�?����H����V9��T�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����d�g�
�
��l�����Ƽ�\��D@��X���u�7�3�f�f�o�(���&�ד�@��Y1�����u�'�6�&��3�%����ѓ�lV�^ �����
�
�
�y�>�����&Ĺ��J��Y1�����b�0�c�u�'�.��������l��h��*���4�
�<�
�$�,�$����ד�@��B�����2�6�0�
��.�N������R��^	������
�!�e�1�0�N�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����I����[��=N��U���u�u�u� ���A����֓�F���'���0�b�0�c�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��E���8�l�|�!�2�}�W���Y���F��B��*��e�0�e�1�w�`��������9��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�(�(܁�O�֓�lV��N�U����;�0�b�2�o�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����d�g�
�
��l�K�������T��h��N���u�u�u�0�$�}�W���Y���F��B��*��e�0�e�1�w�`�U���!����k>��o6��-���������U�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�U��F��g�
�
�
�2�}����Ӗ��P��N����u� �
�
�a�m�����ד�@��Y1�����u�'�6�&��-�������T9��R��!���b�3�8�c�w�%����ǹ��lW��1��Yʴ�
�<�
�&�&��(���H����lW�������6�0�
��$�d����A�ƭ�l��h�����
�!�e�3�:�d�}���Y����]l�N��Uʼ�u�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��PӉ��N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�;�!��-��������lV������1�
� �d�n��E���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��M���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(���P�Ƹ�V�N��U���u�u�7�3�d�l�E߁�&ù��F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�7�3�d�l�E߁�&ù��F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���� 9��^��*ۊ�1�'�&�e�k�}����H����lT��F�X��1�"�!�u�~�W�W���T�Ʈ�U9��X�*���
�1�'�&�f�<����Y����V��C�U���7�3�f�d�e��(ށ�����@W��D�����:�u�u�'�4�.�_���
����@��d:��݊�&�
�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
�ߓ�@��N��*���
�&�$���)�G������F�U�����u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����V����ߊu�u�u�u�w�}����&����l��h�����d�i�u�%�4�3����Oǹ��F�N�����u�|�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�!�0�u�w�}�W���Y����F ��h_�E���d�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���l�3�8�m�~�)����Y���F�N�� ���
�c�e�0�f�<����
�����T�����c�
�}�u�w�}�������9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�`�;���PӒ��]FǻN��U���u�u� �
��k�G���H����A��N�U���6�;�!�9�a��_���Y�ƨ�D��^����u�u�u�9�2�W�W���Y���F��Q1��D��
�
�
�1�%�.�F��YѾ��l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���7�3�f�d�e��(ށ��ƭ�@�������{�x�_�u�w�(�(܁�O�֓�lW��R^�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�d�����@���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�G�������O��_�����u�u�u�u�w�(�(܁�O�֓�lW��R^��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(܁�O�֓�lW��R^��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F���*ي�c�e�0�d�4�l�����Ƽ�\��D@��X���u�7�3�f�f�o�(���&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�*���
�e�u�%�$�:����&����G_��D��Yʴ�
�<�
�&�&��(���I����l_�N�����;�u�u�u�w�4�W���Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ѓ�@��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�f�t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��t�^������F�N��U���7�3�f�d�e��(ށ������T�����2�6�d�_�w�}�W������F�N��U���7�3�f�d�e��(ށ������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y���� 9��^��*ۊ�d�4�&�2�w�/����W���F�U��F��g�
�
�
�f�<����&����\��E�����;��;�0�`�8�F�������T��h��Yʼ�
�4�2�
���[Ϸ�&����V9��R1�U���&�2�6�0��	��������F��h��*���$��
�!�f�;���UӇ��@��T��*���&�l�3�8�o�}��������B9��h��E���8�l�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�e�~�)����Y���F�N�� ���
�c�e�0�f�9�W������]�� 1��B�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��G�����u�u�u�u�w�}�Wϼ��Փ�T��R1�����h�<�
�4�0��(���B���F������}�%�6�;�#�1����H����C9��P1������&�l�3�:�e�^Ϫ���ƹF�N��U��� �
�
�c�g�8�F���Y����]9��Y	��B���f�_�u�u�w�}����Y�έ�l��D�����
�u�u�%�$�:����&����GQ��D��\���=�;�_�u�w�}�W���Y���� 9��^��*ۊ�d�i�u�;��3��������F�N�����u�u�u�u�w�}�Wϼ��Փ�T��R1�����h�w�����/���!����k>��o6��-����w�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z�������P��h��*���u�&�<�;�'�2����Y��ƹF��B��*��e�0�d�"�f�<����&����\��E�����%�6�y�4��4�(�������@��Q��C���-�!�:�1��(�F��&���R��^	������
�!�d�1�0�F������T9��R��!���l�3�8�m�w�-��������`2��C_�����l�_�u�u�2�4�}���Y���Z �F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Dۊ�&�
�e�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����%�6�;�!�;�l�G������\��h��D��
�g�|�u�%�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ց�
����F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Dڊ�&�
�|�|�w�5��ԜY���F�N�����d�g�
�
��8�W������]��[����_�u�u�u�w�1��ԜY���F�N�����d�g�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�"��(��M����A9��G1��*��
�f�i�u�'�>��������N��N����!�u�|�_�w�}����&����l��E��E��u�8�
�`�1��F���	����F��S�����|�_�u�u�z�}����&����l��E��Dʴ�&�2�u�'�4�.�Y��s���Q��1�Mފ�1�'�&�d�6�.���������T��]���&�2�6�0��	���&���� T�V�����&�$��
�#�i����J����F ��h_�A���1�
�0�
�d�j�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�f��.�(��PӒ��]FǻN��U���u�u� �
��e�C�������F������!�9�c�
��}�W�������V�=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�D܁�
����O��_�����u�u�u�u�w�(�(܁�A�ғ�W��D�I��� �
�
�m�c�<��������Q��N��U���0�&�u�u�w�}�W���Yӄ��lU��V�����0�&�u�h�u��}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��Q1��D��
�0�u�&�>�3�������KǻN�� ���
�m�a�6�g�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C]�����f�|�|�!�2�}�W���Y���F��B��*��a�6�e�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����F ��h_�A���e�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���7�3�f�d�o�����
������T��[���_�u�u� ���O����ד�@��Y1�����u�'�6�&��-�������T9��R��!���f�
�&�
�e�}��������B9��h��A���8�f�|�u�w�?����Y���F��QN��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���f�3�8�f�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ғ�@��G��\ʡ�0�u�u�u�w�}�W�������lW��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����J����9��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�U��F��m�
�d�4�$�:�W�������K��N�����f�d�m�
�f�<����&����\��E�����0�
�a�g�w�-��������`2��C]�����f�y�4�
�>�����*���� R��D��F���!�f�d�m��l�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�f��.�(��PӒ��]FǻN��U���u�u� �
��e�C���Y����V��Y����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���J����^9��G�����_�u�u�u�w�}�W���&����R��N�U���f�d�m�
�f�W�W���Y�Ʃ�@�N��U���u�u�7�3�d�l�Oہ�H���>��o6��-���������/���!����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u� �
�
�o�i� ������]F��X�����x�u�u�7�1�n�F��&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�f�3�8�d�q��������V��c1��Fފ�&�
�f�_�w�}����s���F�^��]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�
�&�
�e�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��]��\���=�;�_�u�w�}�W���Y���� 9��Z�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����R��R_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s�����h]��L���0�e�4�1�2�.�W������9��P1�M���u�u�u�:�9�2�G��s���K��B��*��d�0�e�4�3�8����
������T��[���_�u�u� ���N����֓�W��D�����2�
�'�6�m�-����
ۇ��@��T��*���&�b�3�8�a�}��������B9��h��D���8�d�y�4��4�(�������@��Q��M���%�&�2�6�2��#���Hù��^9��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������lT��1��E���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Dڊ�&�
�|�u�?�3�}���Y���F�U��F��f�
�
�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�f�g�d��(߁�����@W�
N��*���&�
�#�a�f�o�Z������\F��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���؁�
����F��R ��U���u�u�u�u�5�;�D��J¹��9��S�����h�4�
�:�$�����I���W��X����n�u�u�u�w�8����Y���F�N�� ���
�l�d�0�g�<����
���D��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u� ���N����֓�VV��D��ʥ�:�0�&�u�z�}�Wϼ��Փ�
U��R1�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���KŹ��^9��G�����u�u�u�u�w�}�Wϼ��Փ�
U��R1����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�Wϼ��Փ�
U��R1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʷ�3�f�g�f���(���Y����T��E�����x�_�u�u�"��(��H����l��h�����%�:�u�u�%�>����	������D�����
��&�b�1�0�A���	����l��F1��*���d�3�8�d�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1����u�0�<�_�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��C���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��PӉ��N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��h��*���u�'�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�g�;���P����[��=N��U���u�u�u� ���N����֓�VW�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u� ���N����֓�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h]��L���0�e�1�u�$�4�Ϯ�����F�=N��U���
�
�l�d�2�m�ށ�
����l��TN����0�&�<�
�6�(��������T��h^����4� �9�:�#�2�(������Z��V �����!�:�
�g�2�i�W���4����_%��C��*���0�c�u�%�$�:����&����GQ��D��Yʴ�
�<�
�&�&��(���H����lW�������6�0�
��$�d����A�ƭ�l��h�����
�!�e�3�:�d�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u� �
��d�F���I����[�S�����;�4��;�%�1�F݁�&����G��DS�X���_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\ʡ�0�u�u�u�w�}�W�������lT��1��E���u�h�}�h�>���������A	��\��*���:�=�'�h�p�z�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���l�3�8�m�~�)����Y���F�N�� ���
�l�d�0�g�9�W��Q����]9��Y��6���'�9�d�
��q�������A�=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�@��������YNךU���u�u�u�u�"��(��H����l��S��E���;��;�4��3����H����J��C����x�|�_�u�w�}�W������F�N��Uʷ�3�f�g�f���(��E����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u� �
�
�n�l��������@��YN�����&�u�x�u�w�?����K����V9��@�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�����UӃ��G��SZ�� ��l�
�g�u�'�.��������l��1����y�4�
�<��.����&����U��B�����2�6�0�
��.�F߁�
����9F����ߊu�u�u�u�1�u�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���H����lW��N��U���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���b�3�8�c�w�3�W���Qۇ��P	��C1��D��h�0�<�6�9�i����M�Г�O���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���I����l_�G�����_�u�u�u�w�}�W���&���� W��h^�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&���� W��h^�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F���*ي�l�d�0�d�6�9����Y����^��1����m�}�u�u�w�2����I��ƓF�C�� ���
�l�d�0�f�<����
�ƭ�@�������{�x�_�u�w�(�(܁�@�ד�lW��S
�����4�&�2�
�%�>�MϮ�������D�����
��&�b�1�0�A���	����l��F1��*���d�3�8�d�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1����u�0�<�_�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y����F ��h\�D���d�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�~�}����s���F�N�����f�g�f�
������
���F��h�����#�a�g�g�z�l��������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�7�3�d�o�Dށ�&¹��W��D_��Hʴ�
�:�&�
�!�i�F��T����\��XN�N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���Ĺ��^9��N�����u�u�u�u�w�}����J����9��1�����&�u�h�4��2�����ғ�T�_�����:�e�n�u�w�}�Wϻ�
��ƹF�N��U��� �
�
�l�f�8�F�������F�L��W�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�(�(܁�@�ד�lW��R^�����;�%�:�0�$�}�Z���Yӄ��lU��]�����6�e�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ߓ�@��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����
9��Z1�\���!�0�u�u�w�}�W���Yӄ��lU��]�����6�e�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���Yӄ��lU��]�����6�e�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�7�3�f�e�n�(���&����R��P �����&�{�x�_�w�}����&����l��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�j����O�ƭ�l��h�����
�!�d�3�:�l�[Ͽ�&����P��h=�����3�8�m�u�'�.��������l��1����_�u�u�0�>�W�W���Y�ƥ�N������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����c�|�:�u��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�G������O��_�����u�u�u�u�w�(�(܁�@�ד�lW��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(܁�@�ד�lW��R_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F���*ي�l�d�0�d�3�}����Ӗ��P��N����u� �
�
�n�l����¹��@��h����%�:�0�&�>���������A	��\��*���<�
�4� �;�2����&�ԓ�lU�^ �����9�:�!�:��o���Y����R��[-�����
�g�0�b�w�-��������`2��CY�����y�4�
�<��.����&����l ��h_�U���&�2�6�0��	��������F��h��*���$��
�!�g�;���s���Q��Yd��U���u�<�u�}�'�>��������lW������6�0�
��$�l�(���&�����YNךU���u�u�u�u�"��(��H����l��S�����;�4��;�%�1�F݁�&��ƹF�N�����u�}�%�6�9�)���������D�����
��&�d��.�(���Y����l�N��U���u�7�3�f�e�n�(���&���F��h#�� ���:�!�:�
�e�8�F�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����f�g�f�
���F��Y����R��[-�����
�g�0�`�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��Q1��G��
�
�
�d�k�}��������\��X��G���b�_�u�u�w�}����s���F�N�����f�g�f�
���F��YѾ��k>��o6��-���������/���!��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�l�d�2�l� ������]F��X�����x�u�u�7�1�n�E��&����D��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�
�$��[ϻ�����WR��B1�L܊�g�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�f�����P�����^ ךU���u�u�3�}��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�F�������F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��B���8�c�u�;�w�2�_ǿ�&����G9��1�Hʰ�<�6�;�a�1��C���	���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�G������O��_�����u�u�u�u�w�(�(܁�@�ד�lW��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(܁�@�ד�lW��R_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F���*ي�e�
�
�
�3�/�������]F��X�����x�u�u�7�1�n�D����֓�W��D�����2�
�'�6�m�-����
ۇ��@��T��*���&�d�
�&��l�W���
����@��d:�����3�8�d�y�6�����
����g9��Z�����f�u�%�&�0�>����-����9��Z1�\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���Q��1�@���e�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Y���F�N��U���
�
�e�
������
���F��h�����#�a�g�g�z�l��������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�n����H���G��d��U���u�u�u�7�1�n�D����֓�W��D�I���%�6�;�!�;�k�(���Y����W	��C��\�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��_��U���;�_�u�u�w�}�W������� V��R1�����0�&�u�h�6�����&����lV�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�g��(߁�����@V�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����J�ӓ�lV��S
����4�&�2�u�%�>���T���F��Q1��F���0�e�4�1�2�.�(�������A	��N�����&�!�%�'�0�o�N������T9��R��!���d�
�&�
�f�}��������B9��h��*���
�y�!�%�d����JŹ��l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���H����^9��G�����_�u�u�u�w�}�W���&����9��1�����&�u�h�!�'�n�(���H����CW�C��U���;�:�e�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�����g�|�!�0�w�}�W���Y�����h]��Eߊ�
�
�1�'�$�l�K�������T9��^��U���u�:�;�:�g�f�W���Y����_��=N��U���u�u�u� ���Gځ�&ù��W��D_��H����n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϼ��Փ�S��h^�����&�<�;�%�8�8����T�����h]��Eߊ�
�
�0�
�$�4��������C��R�����0�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���J����lW�������6�0�
��$�l�(���&���R��^	������
�!�`�1�0�F���Y����V��=N��U���u�3�}�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�o����H���\������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�g�|�:�w�u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fہ�
����O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�~�}����s���F�N�����f�f�`�0�g�>�G��Y����\��h�����n�u�u�u�w�8����Y���F�N�� ���
�e�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}����&����V9��T����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��^�����6�d�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ԓ�@��B�����2�6�0�
��.�D������F�U�����u�u�u�<�w�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����W���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�}����s���F�N�����f�f�`�0�g�>�F��Y����\��h�����n�u�u�u�w�8����Y���F�N�� ���
�e�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}����&����V9��S_�����;�%�:�0�$�}�Z���Yӄ��lU��[��*ڊ�d�4�&�2��/���	����@��U1��F���0�e�$�y�6�����
����g9��\�����d�u�%�&�0�>����-����l ��h\��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�=�;�_�w�}�W���Y�Ʈ�U9��^�����1�u�h�4��2�����ԓ�l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�7�3�d�n�B���I����[��U1��F���0�e�$�n�w�}�W�������9F�N��U���u� �
�
�g��(߁�H���>��o6��-���������/���!����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u� �
�
�g��(߁��ƭ�@�������{�x�_�u�w�(�(܁�Iƹ��9��1�����
�'�6�o�'�2��������F��h�����
�0�1�'�6����I������D�����
��&�d��.�(��Y����P	��1��*���a�%�y�4��4�(�������@��Q��G�ߊu�u�0�<�]�}�W���Y���N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�f�����H�ƭ�WF��CF�����&�!�e�'�6���������9��S�����;�!�9�d�g�t����Q����\��h��*���u�-�!�:�3����Kǹ��O����ߊu�u�u�u�w�}����&����V9��@�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�?����J�ӓ�lV��R_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F���*ي�e�
�
�
�3�/�������]F��X�����x�u�u�7�1�n�D����ד�W��D�����2�
�'�6�m�-����
ۇ��@��T��*���&�d�
�&��l�W���
����@��d:�����3�8�d�y�6�����
����g9��Z�����f�u�%�&�0�>����-����9��Z1�\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���Q��1�@���d�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Y���F�N��U���
�
�e�
������
���F��h�����#�a�g�g�z�l��������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�n����H���G��d��U���u�u�u�7�1�n�D����ד�W��D�I���%�6�;�!�;�k�(���Y����W	��C��\�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��_��U���;�_�u�u�w�}�W������� V��R1�����0�&�u�h�6�����&����lV�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�g��(ށ�����@V�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����J�ӓ�lW��S
����4�&�2�u�%�>���T���F��Q1��F���0�d�4�1�2�.�(�������A	��N�����&�!�%�'�0�o�N������T9��R��!���d�
�&�
�f�}��������B9��h��*���
�y�!�%�d����JŹ��l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���H����^9��G�����_�u�u�u�w�}�W���&����9��1�����&�u�h�!�'�n�(���H����CW�C��U���;�:�e�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�����g�|�!�0�w�}�W���Y�����h]��Eߊ�
�
�1�'�$�l�K�������T9��^��U���u�:�;�:�g�f�W���Y����_��=N��U���u�u�u� ���Gځ�&¹��W��D_��H����n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϼ��Փ�S��h_�����&�<�;�%�8�8����T�����h]��Eߊ�
�
�0�
�$�4��������C��R�����0�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���J����lW�������6�0�
��$�l�(���&���R��^	������
�!�`�1�0�F���Y����V��=N��U���u�3�}�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�o����H���\������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�g�|�:�w�u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fہ�
����O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�~�}����s���F�N�����f�f�`�0�f�>�G��Y����\��h�����n�u�u�u�w�8����Y���F�N�� ���
�e�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}����&����V9��T����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��^�����6�d�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ԓ�@��B�����2�6�0�
��.�D������F�U�����u�u�u�<�w�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����W���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�}����s���F�N�����f�f�`�0�f�>�F��Y����\��h�����n�u�u�u�w�8����Y���F�N�� ���
�e�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}����&����V9��S_�����;�%�:�0�$�}�Z���Yӄ��lU��[��*ۊ�d�4�&�2��/���	����@��U1��F���0�d�$�y�6�����
����g9��\�����d�u�%�&�0�>����-����l ��h\��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�=�;�_�w�}�W���Y�Ʈ�U9��^�����1�u�h�4��2�����ԓ�l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�7�3�d�n�B���H����[��U1��F���0�d�$�n�w�}�W�������9F�N��U���u� �
�
�g��(ށ�H���>��o6��-���������/���!����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u� �
�
�g��(ށ��ƭ�@�������{�x�_�u�w�(�(܁�Iƹ��9��1�����
�'�6�o�'�2��������F��h�����
�0�1�'�6����I������D�����
��&�d��.�(��Y����P	��1��*���a�%�y�4��4�(�������@��Q��G�ߊu�u�0�<�]�}�W���Y���N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�f�����H�ƭ�WF��CF�����&�!�e�'�6���������9��S�����;�!�9�d�g�t����Q����\��h��*���u�-�!�:�3����Kǹ��O����ߊu�u�u�u�w�}����&����V9��@�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�?����J�ӓ�lW��R_��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s�����h]��Eߊ�
�
�1�'�$�m�K���	����@��A\��N�ߊu�u�x�7�1�n�D����ԓ�W��D����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��^�����4�1�0�&��.����	����	F��X��¡�%�'�2�g�n�q��������V��c1��D؊�&�
�d�u�'�.��������l��h��*���!�%�f�
�"�l�Dف�H���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�F݁�
����O��_�����u�u�u�u�w�(�(܁�Iƹ��9��S�����h�!�%�f��(�F��&���K�
�����e�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��G���!�0�u�u�w�}�W���Yӄ��lU��[��*؊�1�'�&�d�k�}��������
V�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�g��(݁�����@W�
N��-��u�u�u�u�2�9���s���V��G�����_�u�u�7�1�n�D����ԓ�VV�
N��*���&�
�:�<��f�}���Y����F ��h]�*���
�0�u�&�>�3�������KǻN�� ���
�e�
�
��8�(�������A	��N�����&�4�
�0�w�-��������`2��C_�����d�y�4�
�>�����*���� 9��Z1����u�0�<�_�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�d�;���P����[��=N��U���u�u�u� ���Gځ�&����F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�7�3�d�n�B���K����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����F ��h]�*���
�d�4�&�0�}����
���l�N�����f�`�0�g�3���������PF��G�����3�
�
�e���(��Y����Z��D��&���!�g�3�8�f�q��������V��c1��F���8�g�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�)����Y���F�N�� ���
�e�
�
��l�K���	����@��A]��E�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��G�����_�u�u�u�w�}�W���&����9��1��U��3�
�
�e���(��s���F�R��U���u�u�u�u�w�?����J�ӓ�lT��N�Uȍ�������/���!����k>��o6��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����J�ӓ�lT��R_�����;�%�:�0�$�}�Z���Yӄ��lU��[��*؊�0�
�&�<�9�-����Y����V��V�����;�'�&�!�g�/��������F9��1��Yʴ�
�<�
�&�&��(���K����lW�������1�
� �d�e��E���	����l��F1��*���
�&�
�|�w�}�������F���]���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ԓ�@��G�����:�}�<�
�2�8�(߁�����V��Q��Lڊ�g�h�4�
�8�.�(���&���R�������!�9�d�e�j�8�����Փ�F9��Z��G���|�!�0�u�w�}�W���Y����F ��h]�*���
�0�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ʈ�U9��^�����"�d�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʷ�3�f�l�e�2�m��������[��Z��D���2�g�m�}�w�}�W������]ǑN��X��� �
�
�d���(���������^	�����0�&�u�x�w�}����J����l��h�����d�4�&�2��/���	����@��G1�����0�
��&�`�;���Y����Z��D��&���!�d�3�8�f�q��������V��c1��L���8�m�u�%�$�:����&����GW��Q��L�ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�6�����
����g9��_�����e�|�!�0�w�}�W���Y�����h]��Dڊ�
�
�1�'�$�l�K���	����@��AX��F��x�d�1�"�#�}�^�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�t����Y���F�N��U���
�
�d�
������
���F��h�����#�a�g�g�z�l��������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�7�3�d�d�G���I����A��N�U���6�;�!�9�a��_���Y�ƨ�D��^����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���N����lP����ߊu�u�u�u�w�}����&����V9��V
�����u�h�4�
�8�.�(���M���K�
�����e�n�u�u�w�}����Y���F�N��U���
�
�d�
������
���F��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�n�N����֓�VV��D��ʥ�:�0�&�u�z�}�Wϼ��Փ�V��h^��ڊ�&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�Eف�
����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���O����lT��G�����_�u�u�u�w�}�W���&����9��1��E��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����J����l��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�� ���
�d�
�
��8�W�������A	��D�X�ߊu�u� �
��l�(���&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�*���
�e�u�%�$�:����&����G_��D��Yʴ�
�<�
�&�&��(���I����l_�N�����;�u�u�u�w�4�W���Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ѓ�@��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�f�t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��t�^������F�N��U���7�3�f�l�g�8�G���H���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U��� �
�
�d���(���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z�������
W��R1�����&�<�;�%�8�8����T�����h]��Dڊ�
�
�d�4�$�:�(�������A	��D�����<�&�a�0�g�}��������l��N��*���;�
�
�
�{�4�(�������V9�������6�0�
��$�j����O�ƭ�l��h�����
�!�d�3�:�l�[Ͽ�&����P��h=�����3�8�m�u�'�.��������l��1����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�e�|�!�2�}�W���Y���F��B��*��
�
�
�d�k�}��������l��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$����������O��_�����u�u�u�u�w�(�(܁�Hù��9��R�����4�;�
�
��f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�m�|�#�8�W���Y���F���*ي�d�
�
�
�f�a�W���>����lR��h\�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�?����@�֓�lV��N�U����<�&�a�2�m�}���Y���V
��d��U���u�u�u�7�1�n�N����֓�F�L��-���������/���!����k>��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�7�1�n�N����֓�VW��D��ʥ�:�0�&�u�z�}�Wϼ��Փ�V��h^��ۊ�&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�@������V��T��A���
�a�c�%�{�<�(���&����l5��D�*���
�e�u�%�$�:����&����G_��D��Yʴ�
�<�
�&�&��(���I����l_�N�����;�u�u�u�w�4�W���Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��^��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�������R��X ��*���
�u�u�-�#�2�ہ�����9��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�l�3�8�o�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��G��\ʡ�0�u�u�u�w�}�W�������l_��h��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W�������
W��R1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N�����l�e�0�d�6�9����Y����^��1����m�}�u�u�w�2����I��ƓF�C�� ���
�d�
�
��9����HӇ��Z��G�����u�x�u�u�5�;�D��I����l��E��D���&�2�
�'�4�g��������C9��P1������&�b�3�:�k�W���
����@��d:�����3�8�d�y�6�����
����g9��1����u�%�&�2�4�8�(���
����U��GךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����W��D��E���!�0�u�u�w�}�W���Yӄ��lU��^��*ۊ�1�'�&�d�k�}��������EP��F�X��1�"�!�u�~�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:�����3�8�l�|�#�8�W���Y���F���*ي�d�
�
�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�f�l�g�8�F�������F������!�9�c�
��}�W�������V�=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�@��������YNךU���u�u�u�u�"��(��&����R��R��U��4�
�:�&��+�C��K�����Y��E��u�u�u�u�2�.�W���Y���F���*ي�d�
�
�
�3�/���E����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�7�3�f�n�m��������@��YN�����&�u�x�u�w�?����@�֓�lW��R^�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�����H���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�E�������O��_�����u�u�u�u�w�(�(܁�Hù��9��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�5�;�D��I����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��B��*��
�
�
�0�w�.����	����@�CךU��� �
�
�d���(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:��݊�&�
�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
�ߓ�@��N��*���
�&�$���)�G������F�U�����u�u�u�<�w�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�|�~�}����s���F�N�����f�l�e�0�f�>�F��Y����\��h�����n�u�u�u�w�8����Y���F�N�� ���
�d�
�
��8�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}����&����V9��S_�����;�%�:�0�$�}�Z���Yӄ��lU��^��*ۊ�d�4�&�2��/���	����@��Y1�����a�0�d�u�9�����M����F��h)�����
�
�y�<��<����&������D�����
��&�b�1�0�A���	����l��F1��*���d�3�8�d�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1����u�0�<�_�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y����F ��hW�*���
�d�i�u�9�����M����l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�m����@����[��=N��U���u�u�u� ���F߁�&¹��Z�^ �����
�
�
�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�����m�|�!�0�w�}�W���Y�����h]��Dڊ�
�
�d�i�w�3�0���
�ғ�lU��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�7�1�n�N����ד�F���2���&�a�0�d�]�}�W���Y����l�N��U���u�7�3�f�n�m�������D��o6��-���������/���!����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�7�3�f�n�m��������@��YN�����&�u�x�u�w�?����@�֓�lW��R_�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�`�;���Y����P	��1��*��c�%�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
�ߓ�@��N��*���
�&�$���)�G������F�U�����u�u�u�<�w�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����V���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9����Q����\��h��*���u�-�!�:�3����@Ź��O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�m�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����
O�N�����u�u�u�u�w�}����J����l��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}����&����V9��@�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��Q1��L���4�1�
�0��(�C���	�����T�����c�
�}�u�w�}�������9F���*ي�`�
�1�'�$�m�K�������l ��[�*��g�x�d�1� �)�W���s���K�U��F��l�4�1�0�$�}����Ӗ��P��N����u� �
�
�b�����
�ד�@��Y1�����u�'�6�&��(�(܁�Lʹ��W��R	��F��u�%�&�2�4�8�(���
�ԓ�@��N��*���
�&�$���)�(���&����C9��P1������&�a�3�:�n�W���
����@��d:��ߊ�&�
�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����l�l�4�1�2�.�W������]��[�*���u�u�u�:�9�2�G��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�`�3�8�c�t����Y���F�N��U���
�
�`�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�f�l�n�<����
�����T�����c�
�}�u�w�}�������9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�;���PӒ��]FǻN��U���u�u� �
��h�(�������Z�U��F��l�4�1�
�2��D��s���F�R��U���u�u�u�u�w�?����@�ߓ�W��D�I����w�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z�������
S��T����2�u�'�6�$�s�Z�ԜY�Ʈ�U9��[�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���HĹ��^9��G�����u�u�u�u�w�}�Wϼ��Փ�_��R^��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(܁�Lʹ��F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���Q��1�L���d�4�&�2�w�/����W���F�U��F��l�6�d�4�$�:�(�������A	��D�����y�4�
�<��.����&����U��B�����2�6�0�
��.�A������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�a�_�w�}����s���F�^��]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�~�2�W���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���O����lS���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�N�����u�u�u�u�w�}����J����l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�"��(��&����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ʈ�U9��[�����&�<�;�%�8�8����T�����h]��@ӊ�d�4�&�2��/���	����@��Y1��*؊�
�y�<�
��o���Y����e9��R1�U����
�
�
�{�<�(���&����l5��D�����d�u�%�&�0�>����-����l ��h[����<�
�&�$���ہ�
������D�����
��&�`�1�0�C�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�a�;���PӒ��]FǻN��U���u�u� �
��h�(��E�ƥ�l6��1��F�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ӓ�@��G�����_�u�u�u�w�}�W���&����
9��R������g�0�g�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��Q1��L���1�u�h�<���E���H���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���7�3�f�l�n�9�W������lT��h^�U���u�u�0�&�w�}�W���Y�����h]��@ӊ�d�i�u����/���!����k>��o6��-������n�w�}�W�������U]�N�����%�:�0�&�]�W�W���Tӄ��lU��W�����&�<�;�%�8�8����T�����h]��@ӊ�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K����lW�R�����`�3�
�a�`�-�[Ͽ�&����P��h=�����3�8�`�u�'�.��������l��h��*���4�
�<�
�$�,�$���ƹ��^9��=N��U���<�_�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�3�8�f�}��������K��X ��*���d�b�
�g�j�<�(���
����9��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���ƹ��^9��G�����u�u�u�u�w�}�Wϼ��Փ�_��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(܁�Lʹ��F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����f(��r����
�
�
� �e�l�(��E��ƹF�N�����
�:�
�:�'�o�(���&����P�������0�
�8�f������O���F�_��U���0�_�u�u�w�}��������Z9��h\�B���n�u�u�0�>�>��������W��N�U��u�=�;�}�e�/���I���R��X ��*���
�|�0�&�w�m�L���YӃ��G��S\�� ��a�
�g�i�w�l�W����Υ�l
��q��9���
�
�0�
�d�d�JϿ�&����G9��1�U���0�w�w�_�w�}��������U��\�����h�w�w�"�2�}�ށ�����^������!�9�f�a�w�1����[���F��^�����3�
�a�c�'�}�J���[ӑ��]F��E�����!�'�
�d������J�����T�����g�g�u�9�2��U�ԜY�Ʃ�Z��Y
�����a�b�%�u�j��Uϩ�����l��h_�@��4�
�:�&��+�(�������V�=N��U���!�:�1�3��l�G���Y���D��_��]���'�2�d�d�w�}��������ET��N�����e�n�u�u�1��2���-����V��Q��E���%�u�h�_�w�}�W���	����@��A]��Eʢ�0�u�!�%�a����J����V�
N��R���9�0�_�u�w�}�W���&����l�N��*����� �
�a�;�(��J����[�N��U���7�3�f�g�d��(ށ�Iӑ��]F��[1��*���
�:�%�f���(���&����V�
N��R���9�0�_�u�w�}�W���&����T��G\�U���3�
�� ������K����lW��1��U��7�3�f�l�g�8�F���B��� ��C��D��g�f�3�
�g�l����D���F�N��*����'��:��j��������U��@��U¡�%�b�
� �e�i�(��I���W����ߊu�u�u�u���;���6����9��P1�G��u�u�3�
�2�0�(��&ǹ��lT�� 1��U��_�u�u�u�w�1��������\�� 1��D���2�g�a�u�?�3�_���&�֓�V��[�E���u�d�|�0�$�}�W���Y����`9��{+��:���`�
�0�
�a�k�}���Y����~3�� ����
�
� �d�c��D��Y���F�������;� �
�c�;�(��H����D��F�����%�
�
� �f�n�(��I���W����ߊu�u�u�u�"��(��&����BV��N�������g��#�e�(���H����CW�
N��'���9�
�a�3��j�N���B��� ��O#��!ػ� �
�a�<��%�(���&����R��G\��Hʦ�1�9�2�6�!�>��������V��h<�� ���&�3�
�c�f�-�^�������]��V�����
�#�m�f���^�ԜY�ƪ�l��{:��:���m�
�;�3��-�(���H����CU�
NךU���u�u�0�
���(�������R��Q��C���%�u�=�;��8�(���K����F9��Y��G��u�u�d�|�2�.�W���Y�����h��*��� �d�d�
�d�W�W����Փ�
S��V
�����u�h�!�%�$�;�(��A����F�N�����u�|�_�u�w�?�D��L����W��D_��Hʡ�%�f�
�0��j�O��T����\��XN�N�ߊu�u�x�3���N�������@��YN�����&�u�x�u�w�;�(܁�@�Փ�VV��D�����:�u�u�'�4�.�_�������C9��P1������&�b�3�:�k�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������9F�N��U���u�7�f�d�b�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����
�l�f�6�g�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�1��(��J������^	�����0�&�u�x�w�}����&����l��h�����%�:�u�u�%�>����	������D�����
��&�f��.�(��s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�e����J�����YNךU���u�u�u�u�5�n�F��&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�3�
�
�n�n���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�;�(܁�@�Փ�F���*ي�m�a�$�n�]�}�W������_��h��U���<�;�%�:�2�.�W��Y����Q9��W�*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&���� Q�N�����;�u�u�u�w�4�W���Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��Y��\���=�;�_�u�w�}�W���Y����lW��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����Q9��^�����4�1�0�&�w�`��������_��F�X��1�"�!�u�~�W�W����Փ�S��h^�����&�d�i�u�:��C�������N��N����!�u�|�_�w�}�Z����Փ�S��h^�����&�<�;�%�8�8����T��� ��1�@���e�6�e�4�$�:�(�������A	��D�����y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h_��\ʡ�0�u�u�u�w�}�W������� V��R1����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�Wϸ�&����9��1��E��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����
�e�
�
��8�W�������A	��D�X�ߊu�u�7�f�d�h�����ד�@��Y1�����u�'�6�&��-�������T9��R��!���f�
�&�
�b�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�c�3�:�n�^�������9F�N��U���u�7�f�f�b�8�G���H���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���7�f�f�`�2�m���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�;�(܁�Iƹ��9��R�����
�c�`�0�g�,�L�ԜY��� ��1�@���e�"�d�4�$�:�W�������K��N�����
�e�
�
��8�(�������A	��N�����&�4�
�0�w�-��������`2��C]�����f�|�u�u�5�:����Y�����F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�f�|�~�}����s���F�N�����
�e�
�
��8�W������]��[����_�u�u�u�w�1��ԜY���F�N��*ي�e�
�
�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�7�d�n�B���H����A��N�U���
� �d�m��l�E��Hӂ��]��G�U���3�
�
�e���(�������Z�C��Fފ�0�
�b�m�e�p�FϺ�����O��=N��U���3�
�
�e���(���Y����T��E�����x�_�u�u�5�n�D����ד�VV��D�����:�u�u�'�4�.�_�������C9��P1������&�g�3�:�l�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������9F�N��U���u�7�f�f�b�8�F���I���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���7�f�f�`�2�l���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϸ�&����9��1��Dʴ�&�2�u�'�4�.�Y��s���U��h]�*���
�0�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��[��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� P��D��@���u�=�;�_�w�}�W���Y�ƪ�lU��[��*ۊ�0�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����lU��h��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN�����f�`�0�d�3�}�Jϲ�&����
S��h_��E�ߠu�u�x�u�5�n�D����ד�VW��D��ʥ�:�0�&�u�z�}�Wϸ�&����9��1��D���&�2�
�'�4�g��������C9��N��*���
�&�$���)�A�������9F����ߊu�u�u�u�1�u�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���O����lU��G�����u�u�u�u�w�}�Wϸ�&����9��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����V9��@�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��h]��Eߊ�
�
�1�'�$�m�K�������lW��1��]���u�u�:�;�8�m�L���YӀ�� 9��1��G���1�0�&�u�j�)���&����Q��\��U���:�;�:�e�l�W�W���TӀ�� 9��1��G���e�4�&�2�w�/����W���F�Q��*��
�
�
�0��.����	����	F��X��´�
�0�u�%�$�:����&����GT��D��\���u�7�2�;�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��D���u�=�;�_�w�}�W���Y�ƪ�lU��[��*؊�0�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����lU��h��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���7�f�f�`�2�o�������]F��X�����x�u�u�3���Gځ�&����9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�c�3�:�n�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�f��.�(��P�Ƹ�V�N��U���u�u�3�
��m�(���&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�3�
�
�g��(݁������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W���J����l��h
�I���!�f�`�l���(��s���K�Q��*��
�
�
�0�w�.����	����@�CךU���7�f�f�`�2�o� �������]9��X��U���6�&�}�%�4�q��������V��c1��F܊�&�
�`�_�w�}����s���F�^��]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�
�&�
�b�t�^Ϫ���ƹF�N��U���7�f�f�`�2�o� ��E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���f�f�`�0�e�*�F��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������U��RN�����u�'�6�&�y�p�}���Y����U��\�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�E܁�
����F��h��*���$��
�!�`�;���UӇ��@��T��*���&�d�
�&��j�W���
����@��d:�����3�8�d�y�6�����
����g9��_�����e�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���L����lT�������6�0�
��$�o�(���&���P
��C1�����:�
�`�0�g�/���I����C9��P1������&�g�
�$��O���	����l��F1��*���e�3�8�g�{�<�(���&����l5��D�*���
�b�u�%�$�:����&����GW��Q��D���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����N��h�����:�<�
�u�w�-��������`2��C\�����g�|�:�u�6�����&����P9��
N��*���
�&�$���)�@�������	�������!�9�2�6�f�`��������V��c1��DҊ�&�
�b�u�%�u��������\��h_��U���&�2�6�0��	���&����_�X�����:�&�
�:�>��W���	����l��F1��*���d�3�8�g�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ԓ�@��G�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��i�W���Q����\��h�����u�u�%�&�0�>����-����9��Z1�\ʺ�u�}�%�6�9�)����I����_9��h(��*���%�f�
�
��8�(��O�ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�b�|�:�w�<�(���
����T��N�����<�
�&�$����������O��EN�����:�&�
�:�>��W���	����l��F1��*���l�3�8�g�~�<����	����@��A_��U���9�9�
�:��2���&����A��X�\���'�}�4�
�8�.�(���&���P
��C1�����:�
�`�0�g�/���I����]�V�����
�:�<�
�w�}��������B9��h��E���8�g�|�|�~�)����Y���F�N����� �d�g�
�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��E�� ��g�
�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�2�%�1��C�������VF��D��U���6�&�{�x�]�}�W���&����T��X�����&�<�;�%�8�}�W�������R��^	������
�!�m�1�0�F������T9��R��!���g�
�&�
�g�}��������B9��h��@���8�g�y�6��)�1���5���� S��h^�����c�c�u�%�$�:����&����GT��Q��G���u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�u�=�9�W�W���Y���F��G1��*��f�:�6�1�w�`��������_��UךU���u�u�9�<�w�u��������_	��T1�Hʴ�
�<�
�&�&��(���H����lT����]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�c�}��������]��[��E��6�
�!��%�����L����l��h\�C���;�u�4�
�8�.�(�������F��h��*���$��
�!�o�;���P���G��d��U���u�u�u�2�'�;�(��J����\��S�����;�!�9�g�g�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��C�������VF�L��W�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�/�(���H����CV��D��ʥ�:�0�&�u�z�}�WϹ�	����R��h�����2�
�'�6�m�-����
۔��lW��B�� ���
�`�
�e�w�-��������`2��C_�����d�y�3�
���8���Lƹ��T9��W����<�
�&�$����������J��G1�����0�
��&�e�����M�ƭ�l��h�����
�!�m�3�:�o�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1�����0�
��&�e�����M�ƣ�N��h�����:�<�
�u�w�-��������`2��C\�����g�|�|�!�2�}�W���Y���F��E�� ��g�
�e�i�w�8�(��O���F�N�����}�4�
�:�$�����&���R��^	������
�!�d�1�0�E���Y����l�N��U���u�2�%�3��i�D���Y����`9��b,�� ���`�'�2�g�c�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�b�~�)����Y���F�N����� �d�g�
�g�a�W���&����
9��d��U���u�0�&�u�w�}�W���Y����A��B1�Gي�e�i�u����/���!����k>��o6��-������n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӁ��l ��Z�*��4�&�2�u�%�>���T���F��G1��*��f�%�
�&�>�3����Y�Ƽ�\��DF����`�y�4�
�>�����*����^��D��B��� �
�
�`�n�,�[ϼ��Փ� U��R1�����4�
�<�
�$�,�$����ד�@��B�� ���
�f�f�0�g�,�[Ͽ�&����P��h=����
�&�
�a�w�-��������`2��C\�����g�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�w�5��ԜY���F�N�����
�a�f�%�w�`����H����9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����M����[��=N��U���u�u�u�'��(�F��&���F��Q1��D��
�
�
�e�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��D���8�g�|�u�?�3�}���Y���F�P�����a�f�%�u�j�?����H����V9��F^�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���A����lW��N�����u�u�u�u�w�}��������U��N�U���
�
�`�l�&�f�W���Y����_��=N��U���u�u�u�'��(�F��&���F��o6��-���������/���!����k>�=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�'�
�"�l�Dށ�IӇ��Z��G�����u�x�u�u�0�-����M�ד�9��D��*���6�o�%�:�2�.��������V��c1��G݊�&�
�c�u�'�.��������l��1����y�3�
������&����S��N��*����g��!�o��(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���KĹ��^9��G�����_�u�u�u�w�}�W���&����U��G^��Hʳ�
����#�h�(���&����l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�i����K���G��d��U���u�u�u�2�'�;�(��H����[��d1�� ���;� �
�a�e�/���N��ƹF�N�����_�u�u�u�w�}�W���&����U��G^��H���������/���!����k>��o6��-���_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������9�������%�:�0�&�w�p�W�������F9��_��D���&�2�
�'�4�g��������V��[�U���&�2�6�0��	���&����P�V�����&�$��
�#�i����K����F ��hW�*���
�e�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�c�~�)����Y���F�N����� �d�f�
�f�a�W���&����9��1��N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ғ�@��G�����u�u�u�u�w�}�WϹ�	����R��h�I���0�
�a�l�]�}�W���Y����l�N��U���u�2�%�3��i�F���Y���k>��o6��-���������/���!����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���2�%�3�
�c�k�����ƭ�@�������{�x�_�u�w�/�(���H����\��S�����;�%�:�u�w�/����Q����Z��D��&���!�d�3�8�d�q����Aù��T9��[����!�%�d�<�%�:�E��Uӕ��l��^��*���
�c�b�u�2����&����T9�� ]����!�%�b�<�%�:�E��UӇ��@��T��*���&�f�
�&��l�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��*���$��
�!�e�;���PӇ��N��h�����#�
�u�u�2����&����T9�� ]�����}�%�6�;�#�1�F��Dӕ��l��Y��*���
�c�l�u�9�}��������]��[��E��&�9�!�%�g�4����K����O�C��U���u�u�u�u�w�:����&����l	��X
��I���%�6�;�!�;�h�C�ԜY���F��D��]���%�6�;�!�;�:���DӇ��@��T��*���&�f�
�&��l�W���Yۇ��P	��C1��D��h�!�%�m��8�(��L�ƭ�WF��G1�����9�d�e�h�$�1����H����V��X�U���u�4�
�:�$��ށ�Y�ƿ�_9��G\�����2�g�c�|�6�9�_�������l
��h^��U���
�8�g�
��8�(��J�ƭ�WF��G1�����9�d�e�h�$�1����N����V��Y�\���=�;�_�u�w�}�W���Y����U��]�����1�u�h�4��2����ƹ��9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�d�����I����[��=N��U���u�u�u�'��(�F��&����W�
N��*���&�
�#�
�l�}�W���YӃ��VFǻN��U���u�u�'�
�"�l�Dف�	����Z�6��-���_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������9�������%�:�0�&�w�p�W�������F9��X��E���&�2�
�'�4�g��������_9��h(��*���%�g�
�
��8�(��O�ƪ�l5��r-�� ���c�'�2�g�e�q��������V��c1��Fۊ�&�
�e�u�"��(��I����l����*���'�2�g�`�{�.����	�ד�l��h\�D���0�
�8�g������O���@��C��L���'�2�g�b�{�.����	�ѓ�l��h\�L���%�&�2�6�2��#���J����^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�>�����*���� T��D��D���;�u�4�
�8�.�(���&���@��C��L���'�2�g�b�~�<����	����@��A_��U���0�
�8�f������O���R��Y��]���6�;�!�9�f�m�Jϭ�����V��h��*��b�|�|�!�2�}�W���Y���F��E�� ��f�
�e�i�w��$���:����lS��E��G��n�u�u�u�w�8����Q�έ�l��D�����
�u�u�%�$�:����&����GU��Q��F���4�1�}�%�4�3����H�����hV�����g�`�|�4�3�u��������EW��S�����8�d�
�
�2��A��Y������T�����d�e�h�&�;�)��������lT�� G�����4�
�:�&��+�(���Y����G��1�����g�b�|�4�3�u��������EW��S�����8�f�
�
�2��A��P�Ƹ�V�N��U���u�u�2�%�1��C���	�����[�����:�%�g�
������L����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!�f�;���P�Ƹ�V�N��U���u�u�2�%�1��C���	�����h]��C���0�d�$�n�w�}�W�������9F�N��U���u�'�
� �f�n�(��E����k>��o6��-���������/���!���9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���'�
� �d�d��FϿ�
����C��R��U���u�u�2�%�1��C���	¹��@��h����%�:�0�&�5�;�D��Kù��9��N��*����'��:��j��������U�������6�0�
��$�n�(���&���G��^�����c�`�u�0��0�Fށ�&����P��N�����%�e�<�'�0�o�A��
����^��h�����c�f�u�0��0�D؁�&����P��N��*���
�&�$���)�E�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�&�2�6�2��#���J����^9��N�����%�6�;�!�;�l�G��
����^��h�����c�f�u�;�w�<�(���
����9��
N�����%�b�<�'�0�o�@�������\�V�����
�#�
�u�w�8�(���Kù��A��X�\���u�=�;�_�w�}�W���Y�ƫ�C9��h_�C���u�h�6�
�#���������l��h��*��b�_�u�u�w�}����Y����C9��Y�����6�d�h�4��4�(�������@��h��*��u�;�u�4��2����¹��F��G1�*���
�c�`�u�9�}��������_��N�����!�%�d�<�%�:�E��PӇ��N��h�����#�
�u�u�2����&����T9��Y�����}�%�6�;�#�1�F��Dӕ��l��W��*���
�c�f�u�9�}��������_��N�����!�%�b�<�%�:�E��P����[��=N��U���u�u�u�'��(�F��&���F��h�����#�g�e�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C]�����f�|�u�=�9�W�W���Y���F��G1��*��c�%�u�h�5�;�D��Kù��9��d��U���u�0�&�u�w�}�W���Y����A��B1�F܊�d�i�u����/���!����k>��o6��-������n�w�}�W�������U]�N�����%�:�0�&�]�}�WϷ�&����\��X��D܊� �d�a�
�e�a�W���&����P9��T��]���<�;�1�<��4�1���5����@9��P1�M���~� �&�2�2�u��������EU��G�U���<�d�3�
�c�n����Dӕ��l
��^�����'� �&�2�2�u�(���&����F�B �����}�%�6�;�#�1�D��P���F��1��*���e�%�u�h�$�9��������G	��B �����}�d�'�2�f�j�^�������]��V�����
�#�
�|�l�}�WϷ�J����W��h�I���!�
�:�<��8��������]��^\�����a�e�u�u�9�4��������]��[��D���_�u�u�
��(�E��&���F��S1�����#�6�:�}�9�4��������T9��_��^ʠ�&�2�0�}�'�>�����ԓ�O��N�����0�0�
�
�2�9����&����
V��N�U��k�;�'�&�#�m�W������K�d��Uʹ�6��d�
�"�l�@ځ�H���U5��y,��1���0�8�g�
�"�l�Aށ�H����F��S�����|�_�u�u�8��(�������U��N�U���4�g�b�
�"�l�@߁�H����W	��C��F��u�u�9�6��l�(���H����CW�
N��#���
�`�3�
�`�m����J�����Y��E��u�u�9�6��l�(���H����CR�
N��#���
�c�3�
�o�h����Iӂ��]��]����u�:�
�
�a�;�(��@����[��h8��G��
� �d�e��l�E���Y�ƨ�D��^����u�:�
�
�`�;�(��L����[��h8��G��
� �d�a��l�D�������T��d��Uʹ�6��d�
�"�l�Bځ�H���C9��[\��B���
�m�d�%��n�Z������\F��d��Uʹ�6��3�
�b�h����DӀ��f(��y*�����
�g�3�
�b�l����Iӂ��]��]����u�!�f�d�o���������F9��1��U��4�
�:�&��+�C��K�����Y��E��_�u�u�x�;��(��A����A��N�����u�'�6�&�y�p�}���Y����lW��1�����&�
�&�<�9�-����Y����V��V�����&�$��
�#�n����J����G9��X�*���'�'�2�g�`�q��������V��c1��D݊�&�
�c�_�w�}����s���F�^��]���6�;�!�9�0�>�F������T9��R��!���f�
�&�
�e�t����Y���F�N��U���f�d�m�
�3�/���E�ƭ�l��D�����g�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�b�1�0�F���Y����l�N��U���u�9�
�
�a�e��������[��C1��D��
�1�'�'�0�o�@��Y���F��[�����u�u�u�u�w�)�D��A˹��W��D^��H����n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϲ�&����^��S
����4�&�2�u�%�>���T���F��h]��C���4�1�0�&��.����	����	F��X��´�
�<�
�&�&��(���J����lU�������6�0�
��$�l�(���&���G��_�����a�d�u�%�$�:����&����GU��Q��F���u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C]�����f�|�u�=�9�W�W���Y���F��h]��C���4�1�0�&�w�`����J¹��T9��_��U���u�:�;�:�g�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�g�~�)����Y���F�N�����d�m�
�1�%�.�F��Y����\��h��A��g�x�d�1� �)�W���s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�b�3�:�l�^������F�N��U���9�
�
�c�o�<����
�����T�����c�
�}�u�w�}�������9F�N��U���0�_�u�u�w�}�W����Փ�^��V
�����u�h�w��l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����G9��X�*���u�&�<�;�'�2����Y��ƹF��C1��D��
�0�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��\����<�
�&�$����������OǻN�����_�u�u�u�w�;�_�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����Փ�@��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��k�^�������9F�N��U���u�!�f�d�o�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����
�c�m�6�g�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�;��(��A������^	�����0�&�u�x�w�}����&����l��h�����%�:�u�u�%�>����	������D�����
��&�f��.�(��Y����Z��D��&���!�b�3�8�f�q��������V��c1��F؊�&�
�d�_�w�}����s���F�^��]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�
�&�
�e�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��X��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�n�^���Y����l�N��U���u�9�
�
�a�e���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���f�d�m�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�!�d�l�Oׁ�H���P
��b ��0���8�g�
�
��(�E��&����9F�C����
�c�m�"�f�<����Y����V��C�U���9�
�
�c�o�*�F���
����C��T�����&�}�%�6�{�<�(���&����l5��D�*���
�d�_�u�w�8��ԜY���F��F��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�t����Y���F�N��U���f�d�m�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�[��*��m�"�d�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�9�
��e�A���I����A��N�����u�'�6�&�y�p�}���Y����lW��1��E���1�0�&�
�$�4��������C��R�����<�
�&�$����������J��G1�����0�
��&�f�����O���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�D܁�
����O��_�����u�u�u�u�w�)�D��MŹ��9��S�����h�4�
�:�$�����K���W��X����n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����Q��D��C���!�0�u�u�w�}�W���Yӊ�� 9��X��*ڊ�1�'�&�e�k�}��������EP��F�X��1�"�!�u�~�W�W���Y�Ʃ�@�N��U���u�u�9�
��e�A���I����A��N�Uȍ�w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���J����9��1�����&�u�&�<�9�-����
���9F���F��a�
�
�
�3�/��������]9��X��U���6�&�}�%�$�:����&����GU��Q��F���4�
�<�
�$�,�$����ѓ�@��B�����d�'�2�g�o�q��������V��c1��GҊ�&�
�b�_�w�}����s���F�^��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�`�t����Y���F�N��U���f�d�a�
������
���F��G1�*���
�a�d�g�z�l��������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�n����J���G��d��U���u�u�u�9���O����֓�W��D�I���%�6�;�!�;�k�(���Y����W	��C��\�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��X��U���;�_�u�u�w�}�W����Փ�R��R1�����0�&�u�h�6�����&����lW�C��U���;�:�e�n�w�}�W�������9F�N��U���u�!�f�d�c��(߁�����@W�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�1�(܁�A�Г�lV��R^�����;�%�:�0�$�}�Z���Yӊ�� 9��X��*ڊ�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���J����^9��N��*���
�&�$���)�@�������9F����ߊu�u�u�u�1�u�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���J����lU��N��U���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�a�t�^Ϫ���ƹF�N��U���!�f�d�a���(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʹ�
�
�m�c�2�m���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϲ�&����P��h^�����&�<�;�%�8�8����T���
��1�A܊�
�
�0�
�$�4��������C��R�����0�u�%�&�0�>����-���� 9��Z1�Yʴ�
�<�
�&�&��(���N����lW�������6�0�
��$�o�(���&���F�U�����u�u�u�<�w�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&���� T���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���b�3�8�d�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ޓ�@�� G��\ʡ�0�u�u�u�w�}�W�������^��h��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W����Փ�R��R1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N��*ي�m�c�0�e�3�}�JϬ�����]ǑN��X���!�f�d�a���(���Y����T��E�����x�_�u�u�#�n�F��&����D��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�m�1�0�E���Y����V��=N��U���u�3�}�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�e����K���F��R ��U���u�u�u�u�;��(��O����l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�#�n�F��&����D��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h]��M���0�d�4�1�2�.�W�������A	��D�X�ߊu�u�!�f�f�i�(���&����V��h�����%�:�u�u�%�>����	����l��F1��*���f�3�8�f�{�<�(���&����l5��D�*���
�c�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�g�~�)����Y���F�N�����d�a�
�
��9����I���R��X ��*���a�g�g�x�f�9� ���Y����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!�`�;���P�Ƹ�V�N��U���u�u�9�
��e�A���H����A��N�U���6�;�!�9�a��_���Y�ƨ�D��^����u�u�u�9�2�W�W���Y���F��h]��M���0�d�4�1�2�.�W��[���9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���!�f�d�a���(���������^	�����0�&�u�x�w�}����&����l��h�����d�4�&�2��/���	����@��G1�����0�
��&�d�����K�ƭ�l��h�����
�!�b�3�:�l�[Ϫ�	����A��Z�Yʴ�
�<�
�&�&��(���A����lT��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h\�\ʡ�0�u�u�u�w�}�W�������^��h��*���'�&�d�i�w�0�(�������^��N�Dʱ�"�!�u�|�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��F���8�f�|�u�?�3�}���Y���F�[��*��c�0�d�4�3�8����DӇ��P	��C1��Cފ�}�u�u�u�8�3���B���F������}�%�6�;�#�1����H����C9��P1������&�d�
�$��A�������9F�N��U���u�!�f�d�c��(ށ�����@W�
N��*���&�
�#�a�f�o�Z������\F��d��U���u�0�&�u�w�}�W���Y����G9��V�*���
�1�'�&�f�a�W͆�[���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����
�m�c�0�f�>�GϿ�
����C��R��U���u�u�9�
��e�A���H����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�f�
�&��o�W���
����@��d:�����3�8�d�|�w�}�������F���]���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�f�3�8�d�t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���!�0�u�u�w�}�W���Yӊ�� 9��X��*ۊ�0�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����lW��1��D���e�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���9�
�
�m�a�8�F���HӇ��Z��G�����u�x�u�u�;��(��O����l��h�����%�:�u�u�%�>����	������D�����
��&�f��.�(��Y����Z��D��&���!�b�3�8�f�q��������V��c1��GҊ�&�
�b�_�w�}����s���F�^��]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�
�&�
�e�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��X��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�m�3�:�o�^���Y����l�N��U���u�9�
�
�o�k�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�!�f�d�c��(ށ������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W���J����9��1��U��'�2�d�`�l�W�W���Tӊ�� 9��X��*ۊ�0�u�&�<�9�-����
���9F���F��a�
�
�
�2���������PF��G�����4�
�0�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF�F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��M���8�g�|�|�w�5��ԜY���F�N��*ي�m�c�0�d� �l�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���F��a�
�
�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�!�d�h�Nځ�&ù��W��D^��Hʡ�%�f�
� �e�n�(��K�����Y��E��u�u�9�
��k�B���I����A��N�U���
�d�'�2�e�e�_���Y�ƨ�D��^����u�x�u�!�d�h�Nځ�&ù��F��D��U���6�&�{�x�]�}�W���J����9��1��E���&�2�
�'�4�g��������C9��N��*���
�&�$���)�B�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&���� R�N�����u�u�u�u�w�}����&����l��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}����L����V9��T�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*ي�c�`�0�e�4�l�����Ƽ�\��D@��X���u�9�
�
�a�h�����ד�@��Y1�����u�'�6�&��-�������T9��R��!���f�
�&�
�f�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�n�^�������9F�N��U���u�!�f�`�n��(߁������T�����2�6�d�_�w�}�W������F�N��U���9�
�
�c�b�8�G���H���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����&����l��h
�I���u�u�u�u�4���������C9��h��*���
�`�c�"�2�}��������l��R	��C��e�u�u�d�~�8����Y���F��R����
�
� �g�o��D�ԶY���F��h]��C���0�e�"�d�6�.��������@H�d��Uʹ�
�
�c�`�2�m� �������]9��X��U���6�&�}�%�4�q��������V��c1��F؊�&�
�d�_�w�}����s���F�^��]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�
�&�
�f�t�^Ϫ���ƹF�N��U���!�f�`�l���(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʹ�
�
�c�`�2�m� ��E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�1�(܁�O�ӓ�lW��S
����i�u�8�
�c�;�(��J����F�N�����u�|�_�u�w�)�D��@ƹ��9��S�����h�!�%�f��8�(��H���W��X����n�_�u�u�z�1�(܁�O�ӓ�lW��R^�����;�%�:�0�$�}�Z���Yӊ�� 9��[��*ۊ�0�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���Jƹ��^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h]�\���=�;�_�u�w�}�W���Y����lS��1��D���e�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������P��h��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���!�f�`�l���(���Y����T��E�����x�_�u�u�#�n�B��&����P��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�g�1�0�D���Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�d�����H���G��d��U���u�u�u�9���A����ד�VW�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�!�d�h�Nځ�&¹��F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����lS��1��D���u�h�3�
���8���Lƹ��T9��W����u�x�9�
��k�B���H������^	�����0�&�u�x�w�}����&����l��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�n�(���&���F�U�����u�u�u�<�w�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&���� W�G�����_�u�u�u�w�}�W���J����9��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����l��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��C1��@��
�
�
�1�%�.�G��Y���� R��B1�Fي�d�g�x�d�3�*����P���F��h]��C���0�g�4�1�2�.�W������9��P1�M���u�u�u�:�9�2�G��s���K��C1��@��
�
�
�0�w�.����	����@�CךU���!�f�`�l���(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�f�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�
�&�
�c�t�W������F�N��Uʹ�
�
�c�`�2�o���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���f�`�l�
������DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���J����9��1��Dʴ�&�2�u�'�4�.�Y��s���_��h[�@���g�6�d�4�$�:�(�������A	��D�����y�4�
�<��.����&����l ��h]����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��Q��F���|�!�0�u�w�}�W���Y����G9��X�*���
�0�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ơ�lU��W�����6�d�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʹ�
�
�c�`�2�o����DӅ��q3��{+�����m�0�g�3��l�D���B���F���F���l�
�
�
�2�}����Ӗ��P��N����u�!�f�`�n��(݁�¹��@��h����%�:�0�&�6�����	����l��F1��*���g�3�8�f�~�}�Wϼ���ƹF�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�n�^���Y����l�N��U���u�9�
�
�a�h�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�!�f�`�n��(݁������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W�������U��Y�����h�w�w�"�2�}����/����U��Z�����u�%�6�;�#�1�O���PӃ��VF�UךU���:�9�&�
�"�l�Nځ�K���V�@��U¹�6��d�
�"�l�Gց�M����C9��Y������|�0�&�w�l�L���Yӈ��_��h��D��
�g�i�u�g�}����Q����e9��h��D��
�a�h�4��2����˹��F��D��D��u�u�;�!�?����L¹��Z�^�����u�9�6��1��B���	���R��X ��*���
��u�9�2��U�ԜY�Ƣ�G��1��*��f�%�u�h�u�� ���Yۊ��l0��1��*��`�%�u�u�'�>��������O��[��W���_�u�u�:�%�.�(���H����CT�
N��Wʢ�0�u�9�6��l�(���H����CW������!�9�g�
�~�8����I��ƹF��X��݊� �d�f�
�e�a�W��Y����N��T1��Dފ� �d�m�
�f�`��������_��h^�����u�e�n�u�w�-�G��&¹��U��Y�����h�_�u�u�w�}��������ET��N�����!�%�`�
�"�l�A؁�K���F�G�����_�u�u�u�w�2�(���K����S��h����u�
�0� �#�j�(���H����CS�
N��&������!�%��E���&����l��_�����:�f�|�s�#�-�Oف�&����V��G]����u�
�0� �#�.����O�ד� F�F��*���&�
�#�e�g�{����/����S��h�N���u�%��9��h����N�֓�F���&�����!�`��8�(��O���F��a��*���3�
�m�`�'�}�Jϼ��Փ�T��R1����u�u�%��;��@���&����l��S�� ���
�c�e�0�f�,�L���YӖ��G��^1��*��g�%�u�h�]�}�W���Y����G9��E1�����d�0�e�'�0�o�O������G��^�����c�`�e�u�w�l�^ϻ�
��ƹF�N��&������!�f�k����I�ޓ� ]ǻN�����
�
�
�
�6�)����&����V��G]��H�ߊu�u�u�u�'�>��������V��@��U¡�%�<�<�<�d����Aƹ��V�
N��R���9�0�_�u�w�}�W�������l
��1�E�ߊu�u�0�
���(���H����CU�
NךU���u�u�%�6�9�)���&������YN�����
�
�
�g�1��B���	����[�I�����u�u�u�u�w�<�(���
����S��^����u�0�
�8�f��(���H����CT�
N�����3�
�l�f�'�}�Ϫ�	����l��X�����3�
�b�l�'�t�}���Y����G��1�����3�
�e�l�'�}�J�������CW��^1��*��l�%�u�:�w�-��������lW�=N��U���
�8�d�
��(�E��&���FǻN��U���9�9�
�:��2���&����A��[�U���;�}�0�
�:�l�(�������W�N��R��u�9�0�_�w�}�W�������l��B1�C؊�f�_�u�u�2����&����^	��V �� ��m�
�g�i�w�)���&����
W��G\��ʦ�9�!�%�d�>�;�(��@����l�N�����%�m�<�3��d�F���Y���@��C��M���1�8�'�4��(�F��&����\��G1�����9�d�d�n�w�}��������l��B1�L݊�g�i�u�!�'�j�(���H����CT��X�����;�!�9�d�f�f�W���
����^��^1��*��d�%�u�h��0�(���&����lW��1��U���u�%�6�;�#�1�F��B�����h��Gڊ�
� �g�e��o�K���
����^��h�� ��l�
�g�4�3�.����	�ߓ�l ��W�*��n�u�u�&�;�)��������V��h�I���u�u�u�u�4���������C9��h��*���
�`�c�"�2�}��������l��R	��C��e�u�u�d�~�8����Y���F��R����
�
� �g�a��D�ԜY�ƿ�_9��G\�����
�e�`�%�w�`�_���&�ߓ�F9��W��Gʴ�1�&�9�!�'�l��������V��h�N���u�&�9�!�'�d����&����l��S�����b�
� �d�a��EϿ�ӕ��l��V��*���g�d�
�g�l�}�Wϭ�����9��Q��C���%�u�h�}�:��D؁�&����U��W�����;�u�0�
�:�l����&����l��d��Uʦ�9�!�%�e�>�;�(��I����[�N��U���6�
�!��%�����H����l��h\�Cʢ�0�u�&�9�#�-�N�������Q��G��U��|�0�&�u�w�}�W���
����^��h�� ��b�
�f�_�w�}��������Z9��h\�B���u�h�}�8��n����@�ߓ�F��SN�����%�m�<�3��d�F���P���F��[1�����<�3�
�e�d�-�W��s���F�V�����
�#�g�b��m�G������@��C��D���'�2�g�c��t�J���^�Ʃ�@�N��U���3�
�0�8��m�(ہ�����9��d��Uʦ�9�!�%�e�>�;�(��I����[�N��U���3�
�0�8��m�(܁�����9�������0�
�8�g������O���F�_��U���0�_�u�u�w�}��������Z9��h\�F���n�u�u�&�;�)��������W��h�I���u�u�u�u�4���������C9��h��*���
�c�b�"�2�}��������l��R	��C��e�u�u�d�~�8����Y���F��R�����
�
� �g�g��D�ԜY�ƿ�_9��GX��*���d�g�
�g�k�}�F������U5��z;��G���!�m�
�;�1�	�������� 9��S�����;�!�9�d��i�G������D��N�����!�%�
�
�"�l�Dށ�K���W�@��U³�
���g��)�Oہ�����J��Q��C���%�u�u�%�4�3����Hƹ��O��[��W���_�u�u�0��0�O������� Q��N�U¦�9�!�%�
��(�F��&����AF��[1��݊�
� �d�f��o�L���Yӕ��l��h�� ��d�
�f�i�w�}�W���YӔ��l��h�� ��l�
�f�"�2�}��������l ��[�*��e�u�u�d�~�8����Y���F��G1�����9�d�
�e�l�}�WϪ�	¹��lW��1��U��}�8�
�g��8��������F9��[��Gʺ�u�8�
�g��8��������F9�� _��G��u�u�!�%�f�j����&����l��S��D���=�;�}�<�9�9����4����])��hV�����-�
�
�
�"�l�Cց�K���@��R
�����;�!�9�d��t�W�������l�N����`�1�8�'�6��(���H����CT�
N�����
�g�<�3��j�@���Y����G��^1��*��� �d�l�
�e�f�W�������Q��R�����<�3�
�m�b�-�W��Q����Z9��h��F���
�m�f�%�w�3�W���&����l��B1�Gӊ�g�n�u�u�#�-�F�������T��^1��*��d�%�u�h��0�(���M����9��h_�L���u�;�u�8���B�������S��G�U���!�%�d�b�>�4����&����l��S��D���=�;�}�:�����Oƹ��[��G1�����9�m��|�2�.�W��B�����h\�����`�f�%�u�j�u��������V��_�����2�d�c�u�8�}��������ET��UךU���8�
�l�3��h�N���Y����G��X	��*���!�'�'�&�-�u��������^��1��*���f�%�|�c�~�f�W�������9��h_�C���u�h�&�1�;�:��������A��M�����;�1�<�
�2��D��U���l�N����
� �d�`��l�K�������T��A�����0�<�0� �$�:����5����u	��{��*���0�
�f�l�{�i�^�ԜY�Ƹ�C9��h��G��
�d�i�u�#�����&����\��R�� �&�2�0�}�e�/���I���O�=N��U���
�`�3�
�f�o����Dӕ��l
��^�����'�'�&�/��3����ۏ��A��Z�\��|�n�u�u�#�-�Bց�����9��R��]���
�
� �d�b��Eϱ�Y����W��^1��*��d�%�|�_�w�}����I����P��h�I���u�u�u�u�6�����&����u ��_��]���
�
� �d�b��E��Y���O��[�����u�u�u�%�4�3����A����F�C��Cۊ� �d�l�
�d�a�W���Y�����hX�����c�d�%�u�?�3�_���&�ߓ�F9��Y��G��u�u�d�|�2�.�W���Y�����hW�����c�l�%�n�w�}����O����lW�� 1��U��}�8�
�
���E���&����l��X�����&�3�
�b�f�-�^�ԜY�Ƹ�C9��h��G��
�g�i�u�#�-�A݁�����P��Y
����� �d�f�
�e�f�W�������9��h_�L���u�h�}�:�%�.�(���H����CT��EN�����`�3�
�m�`�-�^�ԜY�Ƹ�C9��h��D��
�g�i�u�9�)��������W��N��U���9�&�
� �f�d�(��B�����hX�����l�f�%�u�j�u����L����^��h����!�%�c�
�"�l�G؁�K��ƹF��Z��L���
�l�l�%�w�`�_���&�ѓ�F9��]��Gʴ�1�2�%�3��i�A���P���F��G1�*���d�f�
�g�k�}�����ѓ�F9��_��Gʺ�u�:�9�&��(�F��&���9F���*���3�
�l�f�'�}�J�������l ��W�*��4�1�!�%�a����Aʹ��]ǻN�����g�3�
�a�e�2����Y����C9��Y�����g�_�u�u�:��E���&����l��S��&������!�b�����O����F�C��B؊� �d�a�
�f�a�W���&����V��h_��E�ߊu�u�8�
�d�;�(��@����[�C��Bۊ� �d�a�
�e�<�Ϫ�	����U��Z�����_�u�u�8��i����@�ӓ�F�F����
� �d�f��o��������9��h_�B���|�_�u�u�:��B���&����l	��X
��I���%�6�;�!�;�h�E�ԜY�Ƹ�C9��h��D��
�e�i�u���;���6����9��P1�G��u�u�!�%�`����MĹ��Z�U��F��g�
�
�
�g�W�W�������l ��W�*��i�u�!�%�`����Lƹ������*���3�
�a�b�'�t�}���Y����^��B1�A܊�g�i�u�!�'�j�(���&������	��*���d�f�
�g�l�}�WϪ�	����U��[�����1�u�h�4��2����ƹ��9F���*���3�
�a�g�'�}�Jϸ�&����p2��C1�*���
�c�c�_�w�}����@����R��h�I��� �
�
�c�g�8�F���B�����hV�����l�b�%�u�j�u����H����_��h����!�%�b�
�"�l�B݁�K��ƹF��Z��C���3�
�b�d�'�}�J�������l ��X�*��s�%�e�g���(���H����CU�=N��U���
�`�3�
�a�d����DӀ��K+��c\�� ���a�<�
�-���(���H����CT�C��U���;�:�e�n�w�}��������_��N�U���
�:�<�
�2�)�Ǭ�
����F��P ��]���0�
�f�`�{�i�^�ԜY�Ƹ�C9��Q��C���%�u�h�w�u�*����
����WN��h��9����!�m�
�9�8����K����P��h�U���<�;�1�4��2�����ޓ�vO�R��U��n�u�u�!�'�4�݁�&����^��G\��H���w�"�0�u�;�>�!��&����Q��GZ��U���6�;�!�9�o��^ϻ�
���]ǻN�����
�f�<�f��(�F��&���F�N�����9�6��d��(�F��&�����T�����m��|�0�$�}�G��Y����^��h�����
�b�f�%�w�`�U�������
��h8��A���
�b�f�%�w�}��������ET��G�����w�w�_�u�w�0�(���M����9��h_�L���u�h�w�w� �8�Wǲ�����9��h_�@���u�u�%�6�9�)����?����_��^�����u�8�
�
�c�4����A�ߓ�F�L�U���;�}�:�
��k����A�ߓ�F�V�����
�#�f�e�w�1����[���F��G1��ߊ�
� �d�c��o�K���I�ƻ�V�[��#��
� �d�`��l�JϿ�&����G9��]��\ʰ�&�u�d�n�w�}��������lU��Q��@���%�u�h�w�u�*��������lW��Q��@���%�u�u�%�4�3����K������RN��W�ߊu�u�8�
���(���H����CT�
N��Wʢ�0�u�9�6��;�(��L����F��h�����#�
�|�0�$�}�G��Y����^��h��D��
�d�i�u�#�����&����\��R�� �&�2�0�}�%���������W��^1����c�|�c�|�l�8�ϼ�����