-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�?����P��1��@���
�
�c�m�%�0����Y����V��^��U���u�u�u�u�:�0����Y�����^ ��O���7�:�>�n�]�}�W���Y���W��C��U���u�;�0�0�w�`�D��s���F�N�����!�u�u�u�w�3����Y���FǻN��U���u�u�0�
�>�8�W���Y����T��S�����u�n�_�u�w�2����Y���F������u�u�u�;�$�9��������G	��V�����u�:�;�:�g�f�}���Y���F��N��U���o�<�u�!��2���s���F�N��U���u�u�o�:�#�.��������V��EF�����x�u�:�;�8�m�L���Y���F��S
��U���u�u�;�&�3�1��������AN��^
��X���:�;�:�e�l�W�W���Y���P��N��U��<�u�!�
�8�4�L�ԜY���F�S_��U���u�o�<�u�#�����&����\��@����1�"�!�u�~�}�W���Y�����N��U���u�;�&�1�;�:����Y���F��U���u�u�u� �w�)�(�������P��
�����d�1�"�!�w�t�}���Y���F��\N��U���u�u�;�&�3�1����s���]�R �����!�n�_�_�%�5��������G
��QN��3���c�
�
������H����A��^�����;�9�4�1�g�)���
����\��h�����4�<�!�x�w�2����I���@��V�����
�8�u�u�#�����&����\��@����1�"�!�u�~�}����Y����R��NN��U���4�u�e�!�w�8�(������\ ��C
�����
�0�!�'��*����Hӂ��]��G����'�1�#�'�6�1�W���Y�ơ�^9��E����!�<� �0�$�3��������	F��E��N���!�'�7�!�w�$�(���
����	��E��Oʣ�'�4�9�u�$�����&����l��C�� ���'�8�&�,�2�g��������G��U��U���
�!�9�u�1�/�������Q
��^�����,�0�_�!�%�?����(����#��h<��<��������g������ƓQ��YNװ���:�,�4�6�$�����&����A	��D�����e�u�7�2�9�}�W�������l��R�����e�_�x�,�#�8��������R��X��U���u�<�u����9���<�έ�W��P�����<�0�d�u�?�3�W���Y���F��S�����i�u�:�=�%�}�I���^��ƹF����ߊu�u�u�u�w�<�������F��S����u�u�;�u�1�W�Z�������@F��V �����:�_�;�u�%�>���s����^	��h�����e�u�'�6�$�}����Y���T��=N��U���}�9�r�#�9�}�������W������u�u�u�<�w�>�G��^���G��d��U���u�u�u�$�w�`����:����z(��p+�����e�!�%�|�w�}�W���YӃ����=N��U���u�3�_�;�w�/����B���^	��h�����2�4�1�d�w�/����Yۇ��AW�=���ߊu�u�u�1�%�����DӇ��AW��C�����&�&�!�4�$�<�������F��QN��:�������6�9�F���Y����@��_�����_�u�u�u�w�}����H����Z������h�u�e�|�]�}�W������F�N��U���1�'�
�8�w�`����H���F�R ����x�&�;�=�$�.����
����l	��R �����0�&�_�%�:�0��������lW��G�����}�9�|�u�5�:��ԜY�ƥ�N��\I�����4�1�6�>�j�z�P�����ƹF�N�����0�u�u�d�~�)����Y���F�N�����0�u�u�d�~�)����Y���F�N��U���4�}����	�0�������l��G��Hʱ�n�_�u�u�w�}�W����ƥ�l�N��U���u�$�u�h�%�0�4���&����t#��V
��D���%�|�u�u�w�}�Wϻ�ӏ��9F���U���_�;�u�'�4�.�L�Զ����G
��=d�����,���n�"�8�>���W����_	��T1�C���9�n�_�;�>�$����Mà��U9��Q1�����
�c�m�<�]�}�W�������l�N��Uʑ�!��1�=�m��#���+��� T��N��U����1�0�&�6�:�W���7����aF��Z�U���u�u��1�2�.����Y�ƅ�g#��eN�U���_�u�u�:�#�u�W���Y����V��T��;ʆ�����]�}�W���Y����	F��=��*����n�u�u�w�}��������	F��=��*����
��������
����[F�N��"���u�|�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�&�}�W���Y����)��t1��6���}�4�4�<�#�}�W���6����V�=N��U���u�1�'�&�f�g�>���-����t/��a+��:���1�'�&��3�5�Z��=����|F��d��U���u�6�d�o��}�#���6����9F�N��U���u�u�����0���s���F�S_��U���������4���Q����d��_N�Dʑ���u�|�]�}�W���Y���)��=��*����
�����������W��x9��:��|�_�;�u�9�4��Զ����G��B�����u�3�8��c��A���&����_��h_�Mʼ�_�u�u�:�'�3����8����uW��h^��*ߊ�!�`�d�m��<�W���Y���F��X��]���u�u�u�u�w�>���0�Ɵ�w9��p'�����u�u�u�u�w�9����Y����g"��x)��*�����_�u�w�}�W���Y����	F��=��*����n�u�u�w�}�W�������|3��d:��9�������l�}�W���Y�����E_��U���������4���B���F�N��U���u�u�����0���s���F�N�����u������4���:����9F�N��U���u�0�u�u���3���>����F�N��U���$�u�u� �w�	�(���0����p2��UךU���;�u�:�%�9�3�L�Զs����]l�N��3���c�
�
������H����A��bN�U���%�;�;�u��k�G���֓�lS��C1��D��
�4�_�u�w�2�ϳ�	��ƹF�N�����k�6�>�_�w�}�W�������X��S
����_�u�u�u�w�8�W�������F�N�����k�$�y�u�w�}�WϿ����F��S�����u�u�u�u�4�l�J�����ƹF�N��D��u�d�_�u�w�}�W���Y����VW�N��U���$�u�k�$�~�W��������G��B����