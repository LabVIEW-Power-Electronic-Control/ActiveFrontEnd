-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��a��c��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�0�e�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&ù��9��h��U��� �u��
���L���YӖ��l��T�� ����
�����#���Q����\��XN�N���u�%�e�0�f�<�(���Y�ƃ�gF��s1��2���_�u�u�
���W���,�Ɵ�w9��p'��#����u�f�u�8�3���B�����h��*���#�1�o����3���>����F�G1����o������0���/����aF�N�����u�|�_�u�w��(���&����_�!��U���
���n�w�}�������)��=��*����
����u�FϺ�����O��N�����0�a�4�
�;�}�W���Y����)��tUךU���
�
�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���	�֓�lS��G1����������4�ԜY�Ƽ�9��N�:���������4���Y����W	��C��\�ߊu�u�
�
����������f2��c*��:���n�u�u�%�g�8�@��6����g"��x)��*�����}�d�3�*����P���F��1��B���
�9�u�u��}�#���6����9F���*���u�u� �u���8���&����|4�_�����:�e�n�u�w�-�G���A����E
��N��!ʆ�����]�}�W���&����	F��cN��1��������}�D�������V�=N��U���
�
�
�%�!�9�Mϑ�-ӵ��l*��~-�U���%�f�0�e�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����V9��V�����u� �u����>��Y����lU��h_��U���u��
����2���+������Y��E��u�u�%�f�2�l��������|3��d:��9����_�u�u���(���Y����`2��{!��6�����u�f�w�2����I��ƹF��h]��*؊�%�#�1�o��	�$���5����l�N��F���f�o�����;���:����g)��]����!�u�|�_�w�}�(܁�&����l��T�� ����
���l�}�WϮ�J����\��b:��!�����
����_������\F��d��Uʥ�f�0�a�4��1�W���,�Ɵ�w9��p'�����u�
�
�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l��h�����o������0���s���C9��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
���(������)��=��*����n�u�u�'�n���Cө��5��h"��<������}�f�9� ���Y����F�G1�����4�
�9�u�w��W���&����p]ǻN��*ي�
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}�����ޓ�C9��SN�:��������W�W���&����
F��x;��&���������W��Y����G	�UךU���
�
�
�
�'�+���6����g"��x)��N���u�%�f�0�f�}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lU��h_�����9�u�u� �w�	�(���0��ƹF��h]��*��o������0���/����aF�N�����u�|�_�u�w��(���H����E
��N��!ʆ�����]�}�W���&����\��b:��!�����
����_������\F��d��Uʥ�f�0�d�
�'�+���6����g"��x)��N���u�%�f�0�f�}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lU��h_�����9�u�u� �w�	�(���0��ƹF��h]��*��o������0���/����aF�N�����u�|�_�u�w��(���M����E
��N��!ʆ�����]�}�W���&����	F��=��*����n�u�u�6����0�Ɵ�w9��p'�����u�
�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�Ƽ�9��1��*���u�u�����0���s���C9��R1�Oʜ�u��
���f�W���	�ғ�lT��G1�����u��
���L���YӖ��l��T��;ʆ�������8���J�ƨ�D��^����u�
�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�
��}�W���*����|!��d��Uʥ�a�0�a�4��1�W���7ӵ��l*��~-�U���%�a�0�`�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ғ�lS��G1�����u��
���L���YӖ��l��T��;ʆ�����]�}�W���&����R��[
��U��������W�W���&ǹ��F��~ ��!�����
����_������\F��d��Uʥ�a�0�b�4��1�W���7ӵ��l*��~-�U���%�`�0�e�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ӓ�lV��G1�����u��
���L���YӖ��l��T��;ʆ�������8���J�ƨ�D��^����u�
�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�Ƽ�9��1��*���u�u�����0���s���C9��R1�Oʜ�u��
����2���+������Y��E��u�u�%�`�2�n��������z(��c*��:���n�u�u�%�b�8�C��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����h��*���#�1�o��w�	�(���0��ƹF��h[��*���u������4���:����U��S�����|�_�u�u���(ځ�	����\��yN��1�����_�u�w��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�G1�����4�
�9�u�w��$���5����l�N��@���b�o��u���8���&����|4�_�����:�e�n�u�w�-�B���N����E
��N��U���
���n�w�}�������/��d:��9�������w�n�W������]ǻN��*ߊ�
�
�%�#�3�g�>���-����t/��=N��U���
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����R��[
��U��������W�W���&Ź��F��~ ��!�����
����_������\F��d��Uʥ�c�0�e�4��1�W���7ӵ��l*��~-�U���%�c�0�d�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�Г�lW��G1�����u��
���L���YӖ��l��T��;ʆ�������8���Iӂ��]��G�U���%�c�0�g�6�����Y����g"��x)��N���u�%�c�0�d�g�>���-����t/��a+��:���e�1�"�!�w�t�}���Y����V9��V�����u������4�ԜY�Ƽ�9��N�<����
�����#���Q����\��XN�N���u�%�b�0�g�<�(���Y�ƅ�5��h"��<��u�u�%�b�2�l�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����lQ��h_�����1�o��u���8���B�����h��U���������!���6���F��@ ��U���_�u�u�
���(������/��d:��9����_�u�u���(���Y����g"��x)��*�����}�d�3�*����P���F�� 1��F���
�9�u�u���3���>����F�G1����o��u����>���<����N��
�����e�n�u�u�'�j��������WF��~ ��!�����n�u�w�-�@���L����}F��s1��2������u�d�}�������9F���*���
�%�#�1�m��W���&����p]ǻN��*݊�
�u�u����;���:����g)��]����!�u�|�_�w�}�(؁�&Ź��l��T��;ʆ�����]�}�W���&����	F��=��*����
����u�FϺ�����O��N�����0�b�4�
�;�}�W���*����|!��d��Uʥ�b�0�m�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�N����l��A��Oʜ�u��
���f�W���	�ѓ�l_�'��&���������W��Y����G	�UךU���
�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�
�w�}�9ύ�=����z%��N�����0�e�4�
�;�}�W���*����|!��d��Uʥ�l�0�d�o��}�#���6����9F���*���
�%�#�1�m��W���&����p]ǻN��*���0�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}���&����R��[
��U��������W�W���&�֓�lW�'��&���������W��Y����G	�UךU���
�e�0�d�6�����Y����g"��x)��N���u�%�d�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�Ƽ�W��h^�����1�o��u���8���B�����1��D���u��
���(���-��� W��X����n�u�u�%�f��(ށ�	����\��yN��1�����_�u�w��F���K����}F��s1��2������u�d�}�������9F���D���g�4�
�9�w�}�9ύ�=����z%��N����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���H����l��A��Oʜ�u��
���f�W���	����V9��N��U���
���
��	�%���Hӂ��]��G�U���%�d�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�d�2�h�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����lW��R1�����9�u�u����;���:���F��_��*���u������4���:����U��S�����|�_�u�u��l��������WF��~ ��!�����u�n�2�9�}�������V��E�����u�3�8��c��A���Y���F�V�����0���
���6���7����|F��d:��;��u�u�4�!�>�(�ϝ�+����}#��c'��*����:�u�0�6�}�W�������G����U���w��c�e�f�;�Gö�
����V��hZ��=��������`����5����c3��q"��!��������/���I߮��l/��b:��4���-�b�e�e�;�i�C��1����}6��h-��6��`�e�e�e�{��(���,����p.��C��Ɲ�������E���L����.��h=��*���h�f�y����(���D����.��h=��*���h�a�����3���J�ʄ�`9��y1��H��m������#��H�ձ�l�N�����;�u�%�6�9�)�������5��h"��<���h�r�r�_�w�}��������C9��Y�����6�e�o����0���C���]ǻN�����4�!�4�
��.�F������5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�F��Y����\��V ������&�g�3�:�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�n�w�}��������R��c1��F���8�g�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��u�u�6�;�#�3�W���*����9��Z1�Oʆ�������8���K�ƨ�D��^��O���e�e�e�e�g�m�G��I����D��N�����!�;�u�%���ځ�
����	F��s1��2������u�e�}�������	[�^�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���g�u�:�;�8�m�W��[����V��^�E��d�e�e�w�]�}�W���
������d:��݊�&�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����G^��D��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��	��������\��c*��:���
�����l��������\�^�E��e�e�e�d�g�m�G��B�����D��ʴ�
��&�d��.�(���Y����)��t1��6���u�g�u�:�9�2�G���D����V��^�E��e�e�e�e�u�W�W�������]��G1��*���d�3�8�d�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�w�_�u�w�2����Ӈ��`2��C_�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�W�ߊu�u�:�&�6�)����-���� 9��Z1�U����
�����#���Q����\��XN�U��w�e�e�e�g�l�G��I����V�=N��U���&�4�!�4��	���&����U�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I��ƹF��X �����4�
��&�f�����M����g"��x)��*�����}�d�3�*����P���V��^�D��e�e�e�e�g�m�L���YӅ��@��CN��*���&�d�
�&��h�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����W��^�E��e�e�e�n�w�}��������R��c1��D݊�&�
�c�o���;���:����g)��\����!�u�|�o�w�m�G��I����V��^�E��n�u�u�6�9�)����	����@��h��*��o������!���6���F��@ ��U���o�u�e�e�f�m�G��I����V��L�U���6�;�!�;�w�-�$����ߓ�@��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����l�N�����;�u�%���)�G�������	F��s1��2������u�e�}�������	[�^�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�d�1�0�E���Y����)��t1��6���u�g�u�:�9�2�G���D����V��^�E��e�e�e�e�u�W�W�������]��G1��*���g�3�8�g�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y�����d�o�����4���:����V��X����u�h�w�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�d�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�f��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�l�G���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����l'�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h_�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��A]��6��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�d�d�u�W�W�������]��G1�����9�f�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�d�g�l�L���YӅ��@��CN��*���&�
�#�g�d�n�Gۘ�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��_�E��e�e�e�e�g�m�F��I����l�N�����;�u�%�6�9�)���&����S��T��!�����
����_������\F��T��W��d�d�d�d�f�m�F��I����W��^�W�ߊu�u�:�&�6�)��������_��h,��D���g�o�����4���:����U��S�����|�o�u�d�f�l�F��I����V��^�D��e�e�e�n�w�}��������R��X ��*���g�d�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�d�u�W�W�������]��G1�����9�f�
��m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�d�f�m�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Bʱ�"�!�u�|�m�}�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�g�w�2����I����D��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#�b�i�G���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�n�u�u�4�3����Y����\��h��@��e�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����D��N�����!�;�u�%�4�3����A����	F��s1��2������u�`�9� ���Y���F�_�D��n�u�u�6�9�)����	����@��A_��@��o������!���6���F��@ ��U���o�u�e�e�f�l�G��I���9F������!�4�
�:�$�����H���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����d�
�e�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��L�U���6�;�!�;�w�-��������9��N��1��������}�NϺ�����O�
N��E��e�e�e�n�w�}��������R��X ��*���m�f���m��3���>����v%��eN��Bʱ�"�!�u�|�m�}�F��H����W��_�D��u�u�6�;�#�3�W�������l
��1��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�F��H���9F������!�4�
�:�$�����H����g"��x)��*�����}�b�3�*����P���V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g��}���Y����G�������!�9�g�d�m��3���>����v%��eN��U���;�:�e�u�j��F��Y����\��V �����:�&�
�#�e�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B���F��P ��U����
�&�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��w�_�u�u�#�/����Y����V��S��U���!�<�2�_�w�}��������U��R �����u�3�4�
��;���
����_F��L�����_�u�u�<�9�1��������V��c1��D���8�e�o����0���s���@��V�����2�7�1�f�w�}�8���8��ƹF��^	��ʥ�a�0�e�<��4�W���-����t/��=N��U���;�9�%�a�2�m����Y�Ɵ�w9��p'��O���e�n�u�u�$�:����&ǹ��9��h��*���&�2�o����0���s���@��V��*ފ�
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����Z��^	��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u���(ށ����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�a�2�l��������l��T��!�����n�u�w�.����Y����V9��V�����'�2�o����0���C���]ǻN�����9�%�a�0�e�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�i����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��1��*���
�;�&�2�m��3���>����F�D�����
�
�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����V9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�&����V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�<�;�9�'�i��������W9��h��U����
���l�}�Wϭ�����C9��R1�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�c�8�C���&����	F��s1��2���_�u�u�<�9�1�����ғ�A��N��1�����o�u�g�f�W���
����_F��1��A���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��R1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ǹ��9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1�����ӓ�C9��S1��*���u�u��
���L���Yӕ��]��G1�����4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�C���O����@��N��1�����_�u�w�4����	�ғ�lP��E��Oʆ�����m�}�G��Y����Z��[N��A���c�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ف�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9�� 1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ғ�lQ��G1�����
�<�u�u���8���B�����Y�����0�b�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�L����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�h����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��@���d�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ށ�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ӓ�lT��G1�����
�<�u�u���8���B�����Y�����0�g�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�L����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�h����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��@���a�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ہ�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ӓ�lS��G1�����
�<�u�u���8���B�����Y�����0�`�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�L����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�h����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��@���b�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(؁�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ӓ�l^��G1�����
�<�u�u���8���B�����Y�����0�m�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�L����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�h����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��C���e�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(߁�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�Г�lW��G1�����
�<�u�u���8���B�����Y�����0�d�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�N����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�j����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��B���d�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ށ�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ѓ�lT��G1�����
�<�u�u���8���B�����Y�����0�g�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�N����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�j����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��B���a�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ہ�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ѓ�lS��G1�����
�<�u�u���8���B�����Y�����0�`�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�N����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�j����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��B���b�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(؁�	����l��PN�&������o�w�m�L���Yӕ��]��G1�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ѓ�l^��G1�����
�<�u�u���8���B�����Y�����0�m�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�N����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�j����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��N���u�&�2�4�w��(���&����\��c*��:���u�h�r�r�]�}�W�������l_��h^�����1�<�
�<�w�}�#���6����9F������%�l�0�e�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l��h�����o������}���Y����R
��hW��*ۊ�'�2�o����0���C���]ǻN�����9�%�l�0�f�<�(���&����Z�=��*����n�u�u�$�:����&ʹ��9��h��*���2�o�����4��Y���9F������%�d�
�
��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*���0�e�%�0�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�ƿ�T����E���e�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u��m��������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����D���e�<�
�<�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��h��*���2�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�n�w�}�����Ƽ�W��h^�����1�<�
�<�w�}�#���6����9F������%�d�
�
��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�W��h_�����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�H¹��9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1���&����R��[
�����2�o�����4�ԜY�ƿ�T����D���d�4�
�9��/���*����|!��T��R��_�u�u�<�9�1���&����Z��^	��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��l����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
�f�8�E���&����Z��^	��U���
���n�w�}�����Ƽ�W��h\�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
�f�8�D���&����	F��s1��2������u�d�}�������9F������%�d�
�
��/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʥ�d�
�
�
�'�+����&����	F��s1��2���_�u�u�<�9�1���&����R��[
�����o������M���I��ƹF��^	��ʥ�d�
�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����D���a�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����R
��h_�����4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
�f�8�C���&����C��T��!�����u�h�p�z�}���Y����R
��h_�����<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�W��h[�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����l��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�d�
�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����l��h�����o������!���6���F��@ ��U���_�u�u�<�9�1���&����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�<�;�;�-�Fށ�&Ź��l��h�����o������}���Y����R
��h_�����4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�>�(���=����\��B��C���0�e�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�l�}�Wϭ�����T��Q��D܊�g�o�����4���:����U��S�����|�_�u�u�>�3�Ϭ�����\��c*��:���
�����l��������l�N�����u�%�&�2�4�8�(���
�Փ�@��T��!�����n�u�w�.����Y����Z��S
��L���u����l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����I����q)��r/�����u�<�;�9�6�����
����g9��\�����d�o�����4�ԜY�ƿ�T�������7�1�`�a�m��8���7���F��P ��U���
� �b�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��P1�D��������4���Y����W	��C��\�ߊu�u�<�;�;�/���A����g"��x)��*�����}�d�3�*����P���F��P ��U���&�2�6�0��	���&����U�=��*����n�u�u�$�:����	����l��h[�U������n�w�}�����ƫ�C9��1��Dڊ� �c�g�4��2���*����|!��d��Uʦ�2�4�u�'��(�@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʧ�2�b�`�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�m�3�8�`�g�$���5����l�N�����u�%�&�2�5�9�B��CӤ��#��d��Uʦ�2�4�u�'���(���&����_��G1�����u��
���f�W���
����_F��h��*���$��
�!��.�(���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����l5��D�*���
�a�o����0���s���@��V�����2�7�1�`�d�g�5���<����F�D�����'�
�
�
�����@����W	��T��!�����n�u�w�.����Y����Z��D��&���!�l�3�8�f�}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�2�'�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����0�
�l�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��hY�*��o������!���6���F��@ ��U���_�u�u�<�9�1����A���5��h"��<������}�f�9� ���Y����F�D�����'�
� �b�o�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��E��M��o������!���6���F��@ ��U���_�u�u�<�9�1����A���5��h"��<������}�f�9� ���Y����F�D�����%�&�2�6�2��#���Hù��^9��N��1�����_�u�w�4��������T9��S1�F������]�}�W�������C9��P1������&�d�
�$��G��*����|!��d��Uʦ�2�4�u�%�$�:����O���$��{+��N���u�&�2�4�w�8�(��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����<�
�1�
�o�}�W���5����9F������2�%�3�
�e��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��������;� �
�d�h����H����	F��s1��2������u�d�}�������9F������2�%�3�
�d��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������,� �
�e�e�/���I����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
���g��)�E܁�&����V��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��%�"�������U��h��*���b�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�&����P��h=�����3�8�f�o���;���:���F��P ��U���&�2�7�1�`�o�MϜ�6����l�N�����u��-� ��3����J�ғ�F9��X��F��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���5�Ԣ�F��1�����d�d�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����v#��v-�� ���!�f�
�
��8�(��N����g"��x)��*�����}�d�3�*����P���F��P ��U���;�1�
�0�:�.����*����lW��h��*���a�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����l��Z1�������<�d�o�/���J����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
���,�"�����	����l��h_�C��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���5����G9��[�����`�'�2�d�c�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��1���!�g�
�0��h�A��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������
�0�8��%�8����)����A��h��*���g�o�����4���:����U��S�����|�_�u�u�>�3�Ͻ�&����l��Z1�����=�&���$�>�E�������F��d:��9�������w�n�W������]ǻN�����9�3�
�:�2�)��������[��g"�����'�2�d�c�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����P
��X
�����
�4�6�1�3�2����&����T9��V��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�;�3��������R��S�����:�
�
�
�2��B��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����1�
�0�8��.����:����\
��h\�����`�m�o����0���/����aF�N�����u�|�_�u�w�4��������W��R��6���4�0��;�%�1��������^��N��1��������}�D�������V�=N��U���;�9�6�
�8�8����&����R��t�����&�a�'�2�f�e�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��T�����!�'�
�4�4�9��������@9��E��D��u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������G��h-�����1�:�!�:���(���&����\��c*��:���
�����l��������l�N�����u�9�;�1��8����
����W%��C��*���
�0�
�c�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������Y��*���8��&�4�2���������l��h_�M��������4���Y����W	��C��\�ߊu�u�<�;�;�>�(�������^9��D�����;�'�9�&�n�/���H����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʶ�
�:�0�!�%���������]��[1��Dڊ�0�
�c�m�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������_9��S������&�4�0��3����
����A��X�U����
�����#���Q����\��XN�N���u�&�2�4�w����� ����
9��P1�G���u��
����2���+������Y��E��u�u�&�2�6�}��������B9��h��M���8�d�u�u���8���B�����Y�����<�
�1�
�d�}�W���5����9F������3�
����)�A�������F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�B���&����R��C��U����
���l�}�Wϭ�����T��Q1�����3�
�a�
�'�4����Y����)��tUךU���<�;�9�2�'�;�G���L����R��V�����u�u��
���L���Yӕ��]��P�����3�`�3�
�c���������l��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���&����_��Y1�����b�0�d�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��h��*���c�l�<�
�6�:�(؁�&����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�e�3�b�;�(��&����R��hY��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù��9��hX�*����;�0�b�2�i�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �c�n�4�(�������V9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������
9��h<�����
�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����a�
�;��9�8�@���N����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�A�������]��t�����d�
�
�u�w�	�(���0��ƹF��^	��ʲ�%�3�e�3�b�;�(��&����R��[-�����
�g�0�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��h^��*ߊ� �c�l�<��<��������_9��h��U����
���l�}�Wϭ�����T��Q1�����3�
�a�
�9�����:����\
��1��F��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����l ��Z�����4� �9�:�#�2�(������5��h"��<��u�u�&�2�6�}����&ù��9��hX�*����;�4��9�/���&����	F��s1��2������u�d�}�������9F������2�%�3�e�1�h����Mʹ��l+��B�����:�
�g�0�a�g�$���5����l�N�����u�'�
�
���(���O�ߓ�]9��Y��6���'�9�d�
��}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���`�3�
�a��3�0���
�ғ�lV�=��*����
����u�FϺ�����O��N�����4�u�'�
���(ځ�����l��p�����0�d�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h[�� ��l�<�
�4�9��(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�e�3�`�1��Cց�����]��h��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����U��W�����<�&�a�0�c�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���
� �c�l�>�����&ǹ��F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�B���&����Z��V��*ފ�
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�;��<�$�i���Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
�
�
�"�k�N���&����G9��N��1�����_�u�w�4��������lV��h[�� ��l�<�
��e�8�G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���
�
�
� �a�d����/�ԓ�lW�=��*����
����u�FϺ�����O��N�����4�u�'�
���(ځ�����l��g8��*���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����U9��Q��Aӊ�;��
�
��}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���`�3�
�a��3�$���&����	F��s1��2������u�d�}�������9F������2�%�3�e�1�h����Mʹ��l5��1��D��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����l ��Z�����0� �;�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��h^��*ߊ� �c�l�4��8����H����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�A�������G��h\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��(߁�&ƹ��lP��h�����'�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����a�
�%�'�#�/�(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�`�3��i�(�������]9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������
9��h�� ���c�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����l ��h��C���4�
�0� �9�j�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �c�n�<�(�������\��c*��:���
�����l��������l�N�����u�'�
�
���(���O�ߓ�C9��C��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù��9��hX�*���'�!�'�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���
� �c�l�6���������	F��s1��2������u�d�}�������9F������2�%�3�e�1�h����Mʹ��l��N��1�����_�u�w�4��������lV��h_�����l�
�%�&�6�)�Mύ�=����z%��N�����4�u�'�
���(�������9��h���������W�W���������h��*���e�3�
�l��-���� ����g"��x)��N���u�&�2�4�w�/�(���&����l ��W������'�;�0�n�8�G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���
�
�e�3��d�(���)����]��1��D��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����9��hX�*���'�&�!�a�m��3���>����F�D�����'�
�
�
��m����@����l6��P�����0�e�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h_�����l�
�;���<����&����	F��s1��2������u�d�}�������9F������2�%�3�e�1�l�(���O�ԓ�]9��V�����0�e�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h_�����l�
�;��>���������B9��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���I����_��^ ��!���o������!���6���F��@ ��U���_�u�u�<�9�1�����֓�lW��Q��L؊�;��
�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��1��Dڊ� �c�g�4��8����I����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
�g�;�(��&����V��Y1�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-��������U��\�����!�'�
�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��1��Dڊ� �c�g�4��8����J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
�g�;�(��&����VF��d:��9����_�u�u�>�3�Ͽ�&����P��h=����
�&�
�g�m��3���>����F�D�����%�&�2�7�3�d�F��;����r(��N�����4�u�'�
���(ց�����l��D���������W�W���������h��*���
� �b�l�6�����Cӵ��l*��~-�U���&�2�4�u�%��(߁�&ʹ��lQ��h�����,�o�����4�ԜY�ƿ�T��	��*���
�
�
� �`�d����&����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�e�3�n�;�(��&����V��Y1�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-�����ߓ�F9��1��*��� �;�d�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��h��*���b�l�4�
�2�g�$���5����l�N�����u�'�
�
���(���O�ߓ�C9��V�����!�'�
�0�w�}�#���6����	[�I�U���&�2�4�u�%��(߁�&�֓�F9��1��*���'�
�%�&�6�)����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϲ�	����l ��h��B���4�
�!�'��-��������\��c*��:���u�h�r�r�]�}�W�������C9��P1������&�g�
�$��F��*����|!��d��Uʦ�2�4�u�%�$�:����H����	F��x"��;�ߊu�u�<�;�;�:����&����CV�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�j�A���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����<�
�&�$���ځ�
����	F��s1��2���_�u�u�<�9�1��������W9��]��U�����n�u�w�.����Y����Z��D��&���!�c�3�8�f�}�W���&����p]ǻN�����9�4�
�<��9�(��I����|)��v �U���&�2�4�u�'�.��������l��1����u�u��
���L���Yӕ��]��V�����1�
�e�m�m��8���7���F��P ��U���
� �b�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���N�ғ�F��d:��9�������w�n�W������]ǻN�����9�2�%�3��i�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V����� �b�l�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q��@ފ�e�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����S��G^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��%�3�������l ��\�����u��
����2���+������Y��E��u�u�&�2�6�}����&����_��N�&���������W������\F��d��Uʦ�2�4�u�:���N���&����CW�=��*����
����u�EϺ�����O��N�����4�u�8�
���(�������l��N��1��������}�GϺ�����O��N�����4�u�8�
���(���A�Փ�F��d:��9�������w�m��������l�N�����u�0�
�
�����L����	F��s1��2������u�f�}�������9F������!�%�`�<�>�4����O����\��c*��:���
�����}�������9F������&�9�!�%�����L����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�g�>�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʧ�!�g�<�<�>�>��������F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�(���&����l^��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�����&����l_��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�1��:���K����lT��^ �����
�
� �l�d�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��C�����
�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h�� ��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)��������9��T��!�����
����_�������V�=N��U���;�9�!�%�n����J����	F��s1��2������u�`�9� ���Y����F�D�����8�
�l�3��h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��E��
�
�
� �n�j����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����
�
� �l�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����
�a�3�
�`��B��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��������;� �
�d�4�(��� ����F9�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�(���O����F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����l_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��%�"�������U��B1�@���u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������|��Y��*���d�d�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������\��h\�����e�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӊ��l0��1��*��m�%�u�u���8���&����|4�\�����:�e�n�u�w�.����Y���� 9��^1��*���d�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��^1��*���d�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƾ�G9��^1��*���d�a�
�f�m��3���>����v%��eN��Aʱ�"�!�u�|�]�}�W�������^��h��*���3�
�e�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��D���
� �d�b��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1��؊�f�3�
�e�g�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R��*���
�d�
�4�#�>��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�0��0�(�������P��N�&���������W��Y����G	�UךU���<�;�9�%��.����L����V��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�1��:���K����lT��^ �����
�
� �d�g��E��*����|!��h8��!���}�b�1�"�#�}�^�ԜY�ƿ�T����*���3�
�d�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[��ۊ� �d�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��^�� ��g�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����9��h_�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����@Ĺ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Oށ�����9��T��!�����
����_�������V�=N��U���;�9�%�e�g��(�������P��N�&���������W��Y����G	�UךU���<�;�9�!�'�h�(�������R��N�&���������W��Y����G	�UךU���<�;�9�%��.����O����W��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�1��:���K����lT��^ �����0�d�3�
�g�k����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N�����%�
�d�3��l�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�b�<�
�"�l�Oہ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�d�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���-� ��;�"��D�������R��N�&���������W��Y����G	�UךU���<�;�9�2�'�;�(��&����W�=��*����
����u�W������]ǻN�����9�2�%�3��l�(���Cӵ��l*��~-�U���&�2�4�u�'�.��������l��h��*���u��
���f�W���
����_F��h��*���
�a�b�o���2���s���@��V����� �b�g�:�4�9�W���-����t/��a+��:���d�1�"�!�w�t�}���Y����R
��E�� ��g�6�u�u���8���B�����Y�����3�
�g�
�2�g�$���5����l�N�����u�'�
� �`�i����Y����)��tUךU���<�;�9�4������Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����2�7�1�a�d�g�5���<����F�D�����%�&�2�7�3�i�F��;����r(��N�����4�u�%�&�0�?���I����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lR��T��:����n�u�u�$�:����	����l��hZ�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�m�u�u���6��Y����Z��[N��*���
�1�
�e�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��l�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����R��N��:����_�u�u�>�3�Ͽ�&����Q��[�Oʗ����_�w�}����Ӈ��@��U
��D��o�����W�W���������D�����d�l�o����9�ԜY�ƿ�T�������7�1�d�m�m��8���7���F��P ��U���&�2�7�1�f�j�MϜ�6����l�N�����u�%�&�2�5�9�F��CӤ��#��d��Uʦ�2�4�u�%�$�:����K���$��{+��N���u�&�2�4�w�-��������R�,��9���n�u�u�&�0�<�W���
����W��]��U�����n�u�w�.����Y����Z��S
��F���u����l�}�Wϭ�����R��^	�����a�u�u����L���Yӕ��]��V�����1�
�`�u�w��;���B�����Y�����<�
�1�
�b�}�W���5����9F������4�
�<�
�3��A���Y����v'��=N��U���;�9�4�
�>�����N����q)��r/�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��S1�F������]�}�W�������C9��P1����g�o�����}���Y����R
��G1�����1�f�d�o���2���s���@��V�����2�7�1�f�g�g�5���<����F�D�����%�&�2�7�3�n�N��;����r(��N�����4�u�%�&�0�?���A����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lU��T��:����n�u�u�$�:����	����l��h]�U������n�w�}�����ƭ�l��h��*��u�u����f�}���Y����\��CN��3���c�
�
��}�$���YӖ��GF�N��U���4�
�9�u�w��$���5����l�N��Uʴ�
�&�u�u���3���>����F�N�����!�'�u�u���3���>����F�N�����:�0�o����3���>����F�N�����1�0�o����3���>����F�N�����0�1�u�u��}�#���6����9F�N��U����;�0�b�2�m�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y���F��Y1�����b�0�d�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӏ��a��R1����o��u����>���<����N��
�����e�n�u�u�w�}��������9��N�<����
�����#���Q����\��XN�N���u�u�u�<��<����&����	F��=��*����
����u�FϺ�����O��N��U���<�
�4�2���(���Y����g"��x)��*�����}�d�3�*����P���F�N��*���2�
�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���Z��V ��*݊�
�u�u����;���:����g)��]����!�u�|�_�w�}�W�������F��X �����g�0�e�o��}�#���6����9F�N��U����;�4��9�/���&����	F��=��*����
����u�FϺ�����O��N��U���<�
�4� �;�2����&�ԓ�lT�'��&������_�w�}�W�������F��X �����g�0�f�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӏ��~��V�����9�d�
�
�w�}�9ύ�=����z%��N��U���<�
�4� �;�2����&�ԓ�lS�'��&���������W��Y����G	�UךU���u�u�;��9�<�4�������9��N�<����
���l�}�W���Yӏ��~��V�����9�d�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���Z��V��*ފ�
�u�u����;���:����g)��]����!�u�|�_�w�}�W�������]��h��U���������!���6���F��@ ��U���_�u�u�u�w�3�0���
�ғ�lT�'��&���������W��Y����G	�UךU���u�u�;��>�.�C���J����}F��s1��2������u�d�}�������9F�N��U����<�&�a�2�i�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y���F��Y1�����a�0�`�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӏ��t��D1����o��u����>���<����N��
�����e�n�u�u�w�}��������9�� N�<����
�����#���Q����\��XN�N���u�u�u�<��8����Y�ƅ�5��h"��<��u�u�u�u�>��!������/��d:��9�������w�n�W������]ǻN��U���;��
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h>��G���g�o��u���8���&����|4�_�����:�e�n�u�w�}�WϷ�&����l��T��;ʆ�������8���J�ƨ�D��^����u�u�u�;���(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�N������d�0�d�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����C9��C��*���u� �u����>���<����N��
�����e�n�u�u�w�}��������lW�!��U���
���
��	�%���Hӂ��]��G�U���u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�N�����0� �;�f�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���R��R����o������0���/����aF�N�����u�|�_�u�w�}�W�������]9��N��!ʆ�������8���J�ƨ�D��^����u�u�u�%�%�)����Y�ƃ�gF��s1��2������u�d�}�������9F�N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���Y�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�}�WϿ�&����A��T�� ����
�����#���Q����\��XN�N���u�u�u�4��8����H����|3��d:��9�������w�n�W������]ǻN��U���%�'�!�'��l�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���F�V�����u��
���W��Y����]��X�����n�_�u�u�4�0����Ӌ��R��X��E���d�u��u�w�-����s���F�V�����u������4�ԜY���F��h��U���������}���Y���R��C��U���������}���Y���R��X ��Oʚ�������}���Y���R��S��Oʚ�������}���Y���R��R��U��� �u��
���L���Y�����g"�����
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƥ�l6��E�����0�d�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������@��N�<����
���l�}�W���Yӏ��c*��V��*Ҋ�
�u�u����;���:����g)��]����!�u�|�_�w�}�W�������T��D1����o��u����>���<����N��
�����e�n�u�u�w�}��������]9��R1�Oʜ�u��
����2���+������Y��E��u�u�u�u�>���������V��R��@���u��
���(���-��� W��X����n�u�u�u�w�4�(���L����}F��s1��2������u�d�}�������9F�N��U����
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����V��Y1�Oʚ�������!���6���F��@ ��U���_�u�u�u�w�-��������	F��cN��1��������}�D�������V�=N��U���u�%�'�!�%��W���,�Ɵ�w9��p'��#����u�f�u�8�3���B���F������'�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�W���YӇ��P�'��&������|�]�}�W���Y����\��CUװ���u�:�%�;�9�}�6��I����lV��hW��&���u�%�'�u�]�}�W���Y����_�'��&������_�w�}�W���	����\��yN��1�����_�u�w�}�W���
����\��yN��1�����_�u�w�}�W�������	F��cN��1�����_�u�w�}�W�������	F��cN��1�����_�u�w�}�W�������\��b:��!�����n�u�w�}�WϷ�&����	F��=��*����
����u�FϺ�����O��N��U���4�
�0� �9�m�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���F�V�����;�d�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����VF��~ ��!�����u�n�w�}��������]��dװU���6�8�:�0�#�0�1��?�Ъ�9��S
�� ���g�&�f�;��o�D�������CF��=N��U���0�<�u�_�w�}�W���=����}2��r<�U���u�u�����2��0����v4��N��U���1�;�
���}�W���<����9F�N��U���d����m��#���+���F�N�� �����u�u���2���B�����CN��U���u�u�6�>�m��W���&����p]ǻN��U���0�0�u�u���3���>����F�N�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W���H����}F��s1��2������u�d�}�������9F�N��U���:�0�o��w�	�(���0����p2��F����!�u�|�_�w�}�W�������}F��s1��2���_�u�u�u�w�2���6����g"��x)��*�����}�d�3�*����P����F�R �����:�0�!�_�]�}�W���	����GF��qX�3���
�
�4�1�d�3�(���
���� 9��[������u�u�2�9�/����Y���F��sN�<�����_�u�w�}�W���&����vF��~ ��2���_�u�u�u�w�4�G���=���/��r)��N���u�u�u�1�9��>���Y�ƅ�g#��eUךU���u�u�:�!� ��?��0����v4�d��Uʥ�'�u�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�%�.���0�Ɵ�w9��p'�����u�u�u�<�g�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Y�����N�<����
�����#���Q����\��XN�N���u�u�u�6�w�}�9ύ�=����z%��N��U���1� �u�u��}�#���6����e#��x<��F���:�;�:�e�w�f�W�������\��Y��N�ߠu�u�6�8�8�8�ϳ�?����P��1�� ���g�&�f�;��o�D�������CF��=N��U���0�<�u�_�w�}�W���=����}2��r<�U���u�u�����2��0����v4��N��U���1�;�
���}�W���<����9F�N��U���d����m��#���+���F�N�� �����u�u���2���B�����CN��U���u�u�6�>�m��W���&����p]ǻN��U���0�0�u�u���3���>����F�N�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W���H����}F��s1��2������u�d�}�������9F�N��U���o��u����>��Y���F��X��Oʚ�������!���6���F��@ ��U���|�_�u�u�9�}��������9lǻN�����;�;�u��a�m�Fٸ�I����_9��Y��G���f�
�
�4��.�W���Y����V��^�����u�u�u��m��#���+���F�N��8�����o����%�ԜY���F��Y^��<���u�u����f�W���Y����Z��`'��=������]�}�W���Y����l1��c&��U�����u�n�w�}����Y���F�N�����u������4���:����U��S�����|�_�u�u�w�}���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N�����o������0���/����aF�N�����u�|�|�_�w�}��������V��=dװ���;�u�u�2�'�;�G���L����R��N�����0�!�8��c��A���&����F�G��U���u�_�u�u�w�}�������R��[�U���u�u�4�
�$�}�IϿ�&����9F�N��U���&�4�!�h�w�/�(���&����U��W�����4�!�_�u�w�}�W�������X��E��*ڊ�
�
� �c�n�<�(������F�N��*���0�h�u�'���(���&����_��G1�����u�u�u�u�6�����Y����A��h^��*ߊ� �c�l�4��8���Y���F��Y1�����b�0�e�h�w�/�(���&����U��W�����;�0�b�0�g�W�W���Y�ƥ�l4��P��*���u�k�2�%�1�m��������
9��h<�����
�
�y�u�w�}�WϷ�&����V9��R1�H���'�
�
�
�����@����a��R1����_�u�u�u�w�3�%����ѓ�lU�	N�����e�3�`�3��i�(���+����lQ��h]�U���u�u�<�
�6�:�(؁�&�����h��*���
� �c�l�>�����&Ĺ��JǻN��U���;��;�0�`�8�B��Y����U9��Q1�����a�
�;��9�8�@���L���F�N��*���2�
�
�
�w�c�����֓�lS��B1�L���
�4�2�
���[���Y�����e�����0�b�h�u�%��(߁�&ƹ��lP��h��'���0�b�0�b�]�}�W���Y����R��[-�����
�g�0�e�j�}����&ù��9��hX�*����;�4��9�/���&����9F�N��U����;�4��9�/���&����X��E��*ڊ�
�
� �c�n�4�(�������]��[1�*���y�u�u�u�w�4�(�������]��[1�*���u�k�2�%�1�m��������
9��h#�� ���:�!�:�
�e�8�E�ԜY���F��h#�� ���:�!�:�
�e�8�D��Y����U9��Q1�����a�
�;��9�<�4�������9��BךU���u�u�;��9�<�4�������9��N��U���
�
�
�
��(�A�������]��t�����d�
�
�y�w�}�W�������]��t�����d�
�
�u�i�:����I����l ��Z�����4� �9�:�#�2�(�������F�N�����4� �9�:�#�2�(������F��G1��E���`�3�
�a��3�:�������G��h_����_�u�u�u�w�3�:�������G��h_����h�u�'�
���(ځ�����l��z�����;�'�9�d���[���Y�����p�����0�e�h�u�%��(߁�&ƹ��lP��h��2���&�a�0�e�]�}�W���Y����R��hZ��*���k�2�%�3�g�;�B���&����Z��V��*ފ�
�y�u�u�w�}��������9��N��U���
�
�
�
��(�A�������Z��1��G�ߊu�u�u�u�9�����M����[�P�����3�`�3�
�c���������l��d��U���u�<�
�4�9��(���Y����A��h^��*ߊ� �c�l�<��<����&����9F�N��U����<�&�a�2�h�J�������9��1��*��
�;��<�$�i���s���F�^ �����
�
�
�u�i�:����I����l ��Z�����4�;�
�
��q�W���Y����]9��^ ��A���b�h�u�'���(���&����_��Y1�����a�0�b�_�w�}�W�������V��S����3�e�3�`�1��Cց�����V��d��U���u�<�
��e�8�G��Y����U9��Q1�����a�
�;����(��Y���F��Y1��*؊�
�u�k�2�'�;�G���L����R��^ ��#���0�d�_�u�w�}�W���)����V9��
P�����
�
�
�
�"�k�N���&����l��d��U���u�<�
��e�8�D��Y����U9��Q1�����a�
�;����(��Y���F��Y1��*ۊ�
�u�k�2�'�;�G���L����R��^ ��%���0�e�_�u�w�}�W���*����V9��
P�����
�
�
�
�"�k�N���&����l��d��U���u�4�
�0�"�3�G��Y����U9��Q1�����a�
�%�'�#�/�(��Y���F��G1�����
�u�k�2�'�;�G���L����R��V�����;�d�_�u�w�}�W�������]9��
P�����
�
�
�
�"�k�N���&����A��d��U���u�4�
�0�"�3�D��Y����U9��Q1�����a�
�%�'�#�/�(��Y���F��G1�����
�u�k�2�'�;�G���L����R��V�����;�a�_�u�w�}�W�������]9��
P�����
�
�
�
�"�k�N���&����A��d��U���u�4�
�0�"�3�A��Y����U9��Q1�����a�
�%�'�#�/�(��Y���F��G1�����
�u�k�2�'�;�G���L����R��V�����;�b�_�u�w�}�W�������]9��
P�����
�
�
�
�"�k�N���&����A��d��U���u�4�
�0�"�3�N��Y����U9��Q1�����a�
�%�'�#�/�(��Y���F��G1�����
�e�h�u�%��(߁�&ƹ��lP��h�����'�
�e�_�w�}�W���	����F��_��Kʲ�%�3�e�3�b�;�(��&����V��Y1�Y���u�u�u�4��8�J�������9��1��*��
�%�6�|�]�}�WϹ�	����l ��1��*��u�u�:�%�9�3�W���O�֊� ��h��E���u�%�'�u�6�}�}���Y���R��[��Kʴ�
�9�y�u�w�}�WϿ�&����X��G1���ߊu�u�u�u�'�.����D�ƫ�C9��1��Dڊ� �c�g�4��)���Y���F��G1�����k�2�%�3�g�;�F߁�����l��S��Y���u�u�u�4��9���Y����U9��Q1�*���c�g�4�
�3�8�}���Y���R��R��U��2�%�3�e�1�l�(���O�ԓ�C9��V
�����u�u�u�;������&ʹ��F�	��*���
�
�e�3��d�(���)����]��1��E�ߊu�u�u�u�9��;�������V9��
P�����
�
�
�e�1��N݁�����A��R1����_�u�u�u�w�3�������F��G1��E���d�
� �c�e�4�(�������9F�N��U�����4�;���(���GӁ��l ��h��E���
�l�
�;������&˹��JǻN��U���;���4�9��(���Y����A��h^��*���3�
�l�
�9��;�������V9��=N��U���u�;��4�2�3�G���I���T��Q1����
� �c�g�>�����0����V9��=N��U���u�;��<��-����?����S�	N�����e�3�d�
�"�k�E���&����v��T��3���
�`�_�u�w�}�W�������X��E��*ڊ�
�e�3�
�n�����&��ƹF�N�����
�u�k�2�'�;�G���Hù��lP��h��#���y�u�u�u�w�<�(�������[�P�����3�d�
� �a�o��������lV�N��U���4�
�0� �9�l�J�������9��^�� ��g�4�
�0�"�3�F�ԜY���F��h�� ���g�h�u�'���(���I����_��V�����;�g�_�u�w�}�W�������]9��
P�����
�
�
�e�1��N݁�	����F��BךU���u�u�%�6�w�c�����֓�lW��Q��L؊�%�6�|�_�w�}�����֓�l_��B1�L��6�8�:�0�#�0�1��?�Ъ�9��d��Uʥ�'�u�4�u�]�}�W���Y����_�	N��*���y�u�u�u�w�<�(���Y����C9��CBךU���u�u�%�&�6�)�J�������9��1��*��
�%�&�4�#�W�W���Y�ƭ�l��RN��U���
�
�
�
��(�@�������]�N��U���4�
�1�0�j�}����&ù��
9��hY�*���<�9�y�u�w�}�WϿ�&����JF�	��*���
�
�
� �`�d��������9F�N��U���-�e�h�u�%��(߁�&ʹ��lQ��h����_�u�u�u�w�-��������X��E��*ڊ�
�
� �b�n�<�(�������l�N��Uʴ�
�0� �;�f�`�W���&����U9��Q��Eӊ�%�'�!�'��q�W���Y����C9��S����3�e�3�l�1��Gց�	����lǻN��*ڊ�4�1�&�7�d�3�(���
���� 9��[�����c�u�u�:�'�3����8����uW��h^�����&�7�f�;��o���&����_
��DךU���0�0�<�u�6�}�}���Y���z"�	N����u�u�u� ��	�0���G����F�N�����
���u�i�n�[���Y�����1��1���h�u�g�_�w�}�W�������z"��S�F���u�u�%�'�w�<�W�ԜY���F��\N��U���6�>�_�u�w�}�W��������E�����u�u�u�<�g�`�W���&����P��BךU���u�u�<�d�j�}��������l��=N��U���u�%�:�0�j�}��������l	��X
�����u�u�u�0�j�}��������l��=N��U���u�:�!�h�w�/�(���N�Г�O��=N��U���
�4�1�&�5�n����K����9��Q��*���
�c�u�u�8�-����Y����V����*���1�&�7�f�9��E���J����U��h
�����u�0�0�<�w�<�W�ԜY���F��S�D�ߊu�u�u�u���#���Y���l�N��Uʱ�;�
���w�c�D��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��|�u�u�%�%�}����s���F�T��H���%�6�>�_�w�}�W�������X��G1���ߊu�u�u�u�>�m�J�������lQ��h����u�u�u�<�f�`�W���&����T��BךU���u�u�%�:�2�`�W���&����T��G���ߊu�u�u�u�2�`�W���&����T��RBךU���u�u�:�!�j�}��������l��dךU���
�
�4�1�d�3�(���
���� 9��[�����c�u�u�:�'�3����8����uW��h^�����f�;�
�g�$�n�(܁�����@ǻN�����<�u�4�u�]�}�W���Y���F��=N��U���u� �
���}�I��s���F�S��*����u�k�f�{�}�W���Yӂ��9��s:��H���g�_�u�u�w�}����.����[�\��U���%�'�u�4�w�W�W���Y�Ư�XF������_�u�u�u�w�8����GӇ��A��=N��U���u�<�e�h�w��F���H����@��=N��U���u�<�d�h�w��F���K����@��=N��U���u�0�h�u�%����A����9F�N��U���!�h�u�'��(�@���	����9F���*���7�f�;�
�e�.�D݁�&����l��h;�U���:�%�;�;�w��A���Hŀ��l ��U1����g�&�f�
��(����	�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�d�W�W���Y�ƨ�]V��~*��U��f�y�u�u�w�}����&����{F�]����u�u�u�:�#�
�3���D����l�N�����4�u�_�u�w�}�W���Y����C9��\BךU���u�u�0�0�w�c����
��ƹF�N����h�u�
�d�2�l������ƹF�N����h�u�
�d�2�o������ƹF�N����u�'�
� �`�i���Y���F��X��H���'�
� �b�c�-�^�ԶY����lV��Z��Fػ�
�g�&�f������
����F��T�����!�8��a��k�(߁�������\��*���d�8�-�1�'�}�WϹ�������FךU���u�u��h�w�q�W���Y����f+��c/��U��d�_�u�u�w�}����.����[�\�U���u�u�1�;���#���G����9F�N��U���!����j�}�E�ԜY�Ƽ�A��V�����u�u�u�<�g�`�W���&����R��BךU���u�u�<�d�j�}��������l��=N��U���u�:�!�h�w�/�(���N�ғ�O��=N��U���
�8�9�f�9��E���J����^��S�� ��o�6�8�:�2�)����Mà��U9��Q��*���&�f�;�
�e�l������ƹF��R �����4�u�_�u�w�}�W���D����9F�N��U���
���u�i�l�}���Y���W��h9��!���k�f�y�u�w�}�WϺ�¹��w2��
P��G�ߊu�u�u�u�8�)� ���1��� T�N�����u�4�u�_�w�}�W������F��G1��*��
�e�_�u�w�}�W���H���T��Q��Aӊ�d�_�u�u�w�}����D�ƫ�C9��hY�*��n�_�u�u������J���� T��h]��D���-�1�%� �`�g����������Z��Dܳ�e�3� �
�e�.�Dݰ�&�ԓ�l��h
�����u�0�0�<�w�<�W�ԜY���F��S�D�ߊu�u�u�u���#���Y���l�N��Uʱ�;�
���w�c�D��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��|�u�u�%�%�}����s���F�S��U��2�%�3�
�b��G�ԜY���F��Y_��Kʳ�
�:�0�!�%�����
����Z9��1����f�y�u�u�w�}����Y����A��B1�A���|�_�u�u�1�m����&�Ԣ�lU��D1�*ۊ�4�
�&�
�a�}�W���	����GF��qX�3���
�
�8�9�d�3�(���
����9��O1�����u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���g�_�u�u�8�)����Q���F�
��E��u�'�
� �`�e���Y���F��^ �H����;�1�
�2�0��������E��Y�����`�a�_�u�w�}�W������T��Q��@Ҋ�g�n�_�_�]�}�W������F��Y�����u�4�
��1�0�W�������G�������{�x�_�u�w�-�4���
����@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ��U���u�u�u�u�w�}�W�������l ��R������3�8�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����
�
�
�e�1��N݁�	����A��G1�����'�2�4�&�0�}����
���l�N�����e�3�d�
�"�k�E���&����G9��h�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}����&ù��V��B1�G���
�!�'�
�'�.�������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���J����lW��G�����_�u�u�u�w�}�W���Y���T��Q1����
� �c�g�6�����&����G��h��U��4�
�:�&��2����B���F�N��U���u�9�<�u��-��������Z��S�����
�
�
�e�1��N݁�	����W����ߊu�u�u�u�w�}�W���Y�ƫ�C9��1��Dڊ� �c�g�4��)����	����A��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�2�%�1�m��������
9��h�����%�&�4�!�%�:�����Ƽ�\��D@��X���u�2�%�3�g�;�B���&����R��C��*���&�4�!�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӁ��l ��h��*���c�l�4�
�#�/�(���
����l��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����R��D��F���;�u�:�}�6�����&����P9��
N�����e�3�d�
�"�k�E���&����O����ߊu�u�u�u�w�}�W���Y�ƫ�C9��1��@���
�a�
�%�$�<����&����G9��PN�U���6�;�!�9�0�>�F�ԜY���F�N��Uʰ�&�3�}�4��2��������F�P�����3�`�3�
�c����������YNךU���u�u�u�u�w�}�W�������9��1��*��
�%�&�4�#�<�(�������TF������!�9�2�6�g�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���'�
�
�
�����@����@��C1��*���'�
�0�u�$�4�Ϯ�����F�=N��U���
�
�
�
��(�@�������R��V�����
�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����U9��Q��Eӊ�%�&�4�!�6�����&����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���N����lP�N�����u�u�u�u�w�}�W���Y����A��h^��*ӊ� �b�l�4��)����	����A��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���9�<�u�}�'�>��������lW�	��*���
�
�
� �`�d��������F��R ��U���u�u�u�u�w�}�W�������lV��hW�� ��l�4�
�!�%���������V�
N��*���&�
�:�<��f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�d�
�
��-����	����R��P �����&�{�x�_�w�}�(����֓�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u��m��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���K����lT��N�����u�u�u�u�w�}�W���Y���F��h_�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�d�~�)����Y���F�N��U���u�u�u�u��m��������W9��R	��Hʥ�d�
�
�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�d�
�
�
�%�:�����Ƽ�\��D@��X���u�%�d�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h_�����%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u��m��������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�V��h^�����i�u�
�e�2�m�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�d�0�g�<�(���&������^	�����0�&�u�x�w�}���&����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�l�(���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���K����^9��G�����_�u�u�u�w�}�W���Y���F�G1�*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�a�f�}����s���F�N��U���u�u�u�u�'�l�(���&����_��E��I���
�d�0�e�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�d�0�e�'�8�W�������A	��D�X�ߊu�u�
�d�2�m����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1�*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�l�(���&����_�N�����u�u�u�u�w�}�W���Y����lW��R1�����u�h�%�d���L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�d�
����������TF��D��U���6�&�{�x�]�}�W���H����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��F���H����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ԓ�@��G�����u�u�u�u�w�}�W���Y���F���D���d�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�c�t����Y���F�N��U���u�u�u�u�w��F���H����E
��G��U��%�d�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�d�
�
��/�Ͽ�
����C��R��U���u�u�%�d���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���D���d�%�0�u�j�<�(���
���� T��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��F���H����E
��G�����_�u�u�u�w�}�W���Y���C9��h��*���2�i�u�
�f�8�F�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�d�2�o��������V��D��ʥ�:�0�&�u�z�}�WϮ�H¹��9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�Fށ�&����l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��_��U���;�_�u�u�w�}�W���Y���F�N��Dۊ�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W���Y���F��D��]���&�2�7�1�c�d�W������F�N��U���u�u�u�u�w�-�Fށ�&����l��h����u�
�d�0�e�<�(���B���F�N��U���u�u�u�;�w�;�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�d�0�e�-����
������T��[���_�u�u�
�f�8�E�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��Dۊ�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�Fށ�&����l��G�����u�u�u�u�w�}�W���Y�����1��G���0�u�h�%�f��(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�d���(�������A��V�����'�6�&�{�z�W�W���&�ד�lU��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(����Փ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h\�\ʡ�0�u�u�u�w�}�W���Y���F�N��*���0�f�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��h�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(����Փ�C9��S1�����h�%�d�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�d�
����������]F��X�����x�u�u�%�f��(܁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*���0�f�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(����Փ�C9��SG��U���;�_�u�u�w�}�W���Y���F��_��*ي�'�2�i�u��l���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
�f�8�C���&����C�������%�:�0�&�w�p�W���	����V9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}���&����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���F�N����
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�i�@������F�N��U���u�u�u�u�w�}���&����R��[
�����i�u�
�d�2�i������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�d�2�i����Y����T��E�����x�_�u�u��l����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N����
�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`���&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h_�����%�0�u�h�'�l�(���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�f��(ځ�	����l��PN�����u�'�6�&�y�p�}���Y����l��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���H����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���!�0�u�u�w�}�W���Y���F�N��U���d�0�`�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��@�������9F�N��U���u�u�u�u�w�}�W���H����l��A�����u�h�%�d���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�d���(���Ӈ��Z��G�����u�x�u�u�'�l�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���d�0�`�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���H����l��A��\���=�;�_�u�w�}�W���Y���F�G1�*���
�'�2�i�w��F���L���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u��l��������W9��R	�����;�%�:�0�$�}�Z���YӖ��9��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�H¹��9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���u�=�;�_�w�}�W���Y���F�N��Uʥ�d�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�C��Y����l�N��U���u�u�u�u�w�}�WϮ�H¹��9��h��*���2�i�u�
�f�8�A���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
�f�8�A����ƭ�@�������{�x�_�u�w��F���O����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�d�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�H¹��9��h��\���!�0�u�u�w�}�W���Y���F���D���c�%�0�u�j�-�Fށ�&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�i��������W9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���F�N�����0�e�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��m�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ہ�&ù��l��h����u�
�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�a�0�e�'�8�W�������A	��D�X�ߊu�u�
�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hZ��*ڊ�'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���&ǹ��9��h��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������O�C��U���u�u�u�u�w�}�W���YӖ��l��h����u�
�
�
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�a�0�d�4��1�(���Ӈ��Z��G�����u�x�u�u�'�i��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�}�'�>��������lW������6�0�
��$�o�(���&�����YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����d�|�!�0�w�}�W���Y���F�N��U���u�
�
�
��-����	����[��hZ��*ۊ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1��D���0�u�&�<�9�-����
���9F���*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�M����l��PN�U���6�;�!�9�d��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����0�d�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u���(ށ����F��1��D�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lR��h\�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�
�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���g�3�8�g�~�}����s���F�N��U���u�u�u�u�'�i��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����T�����ߊu�u�u�u�w�}�W���Y���F��1��G���
�9�
�'�0�a�W���&����R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����ԓ�A��V�����'�6�&�{�z�W�W���&ǹ��9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
������E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�
�'�0�a�W���&����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�C���J����E
��G��U���<�;�%�:�2�.�W��Y����lR��h]�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ǹ�� 9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GT��Q��G���u�=�;�_�w�}�W���Y���F�N��Uʥ�a�0�f�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��D�������9F�N��U���u�u�u�u�w�}�W���&����R��[
�����i�u�
�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�a�0�d�-����
������T��[���_�u�u�
���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�i��������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�9��1�����h�%�a�0�d�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�a�2�i��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�E�������F��R ��U���u�u�u�u�w�}�W���Y����lR��hZ�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����d�g�u�=�9�W�W���Y���F�N��U���u�%�a�0�c�<�(���&����Z�G1�����4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hZ��*ފ�'�2�4�&�0�}����
���l�N��A���a�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ǹ��9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�a�0�a�4��1�^�������9F�N��U���u�u�u�u�w��(���&����Z�G1����_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h��*���#�1�%�0�w�.����	����@�CךU���
�
�
�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��A���`�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�e�t�W������F�N��U���u�u�u�u�w�-�C���L����E
��G��U��4�
�:�&��2����B���F�N��U���u�u�u�9�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1�����4�
�9�
�%�:�K���&ǹ��9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�M����l��PN�����u�'�6�&�y�p�}���Y����V9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
���(������R��X ��*���g�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lR��h[�����1�|�u�=�9�W�W���Y���F�N��Uʥ�a�0�`�%�2�}�JϮ�M����l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ہ�&Ź��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��R1�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ғ�lP��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�F��Y����l�N��U���u�u�u�u�w�}�WϮ�M����l��A�����u�h�%�a�2�k������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
����������]F��X�����x�u�u�%�c�8�A�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��A���c�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�C���O����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�a�2�k�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(ہ�&Ĺ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�c�8�@���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�d�l�u�?�3�}���Y���F�N��U���u�u�%�a�2�j��������V�
N��A���b�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�b�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�C���N����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1��E���
�9�
�'�0�<����Y����V��C�U���%�`�0�e�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ځ�&ù��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W�� V�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ӓ�lV��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ƹ��9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�8�G��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&ƹ��]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����ד�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�`�0�d�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ƹ��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`�2�l����Y����T��E�����x�_�u�u���(ށ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�B���H����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�`�2�l�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(ځ�&����l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�8�E���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�d�c�u�?�3�}���Y���F�N��U���u�u�%�`�2�o��������V�
N��@���g�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�g�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�B���K����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1��F���
�9�
�'�0�<����Y����V��C�U���%�`�0�f�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ځ�&����l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��[�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ӓ�lU��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ƹ�� 9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�8�D��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&ƹ�� ]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����ғ�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�`�0�a�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ƹ��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`�2�i����Y����T��E�����x�_�u�u���(ہ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�B���M����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�`�2�i�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(ځ�&ƹ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�8�B���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�g�f�u�?�3�}���Y���F�N��U���u�u�%�`�2�h��������V�
N��@���`�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�`�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�B���L����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1��C���
�9�
�'�0�<����Y����V��C�U���%�`�0�c�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ځ�&Ź��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��\�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ӓ�lP��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ƹ��9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�8�A��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&ƹ��]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����ѓ�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�`�0�b�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ƹ��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`�2�j����Y����T��E�����x�_�u�u���(؁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�B���N����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�`�2�j�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(ځ�&˹��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�8�O���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�g�e�u�?�3�}���Y���F�N��U���u�u�%�`�2�e��������V�
N��@���m�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�m�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�B���A����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1��L���
�9�
�'�0�<����Y����V��C�U���%�`�0�l�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ځ�&ʹ��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��W�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ӓ�l_��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ƹ��
9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�8�N��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&ƹ��
]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����֓�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�c�0�e�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ź��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�c�2�m����Y����T��E�����x�_�u�u���(߁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*܊�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�A���I����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�c�2�m�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(ف�&¹��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�a�8�F���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�g�b�u�?�3�}���Y���F�N��U���u�u�%�c�2�l��������V�
N��C���d�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�d�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�A���H����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��E���
�9�
�'�0�<����Y����V��C�U���%�b�0�e�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&ù��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��[�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ѓ�lV��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�8�G��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&Ĺ��]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����ד�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�b�0�d�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b�2�l����Y����T��E�����x�_�u�u���(ށ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@���H����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�b�2�l�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(؁�&����l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�8�E���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�f�f�u�?�3�}���Y���F�N��U���u�u�%�b�2�o��������V�
N��B���g�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�g�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�@���K����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��F���
�9�
�'�0�<����Y����V��C�U���%�b�0�f�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&����l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��\�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ѓ�lU��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ�� 9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�8�D��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&Ĺ�� ]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����ғ�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�b�0�a�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b�2�i����Y����T��E�����x�_�u�u���(ہ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@���M����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�b�2�i�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(؁�&ƹ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�8�B���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�f�e�u�?�3�}���Y���F�N��U���u�u�%�b�2�h��������V�
N��B���`�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�`�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�@���L����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��C���
�9�
�'�0�<����Y����V��C�U���%�b�0�c�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&Ź��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��W�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ѓ�lP��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�8�A��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&Ĺ��]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����ѓ�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�b�0�b�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b�2�j����Y����T��E�����x�_�u�u���(؁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@���N����E
��G�����_�u�u�u�w�}�W���Y���C9��R1�����u�h�%�b�2�j�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
��-����	����R��P �����&�{�x�_�w�}�(؁�&˹��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�8�O���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$����������O�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�f�b�u�?�3�}���Y���F�N��U���u�u�%�b�2�e��������V�
N��B���m�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N�����0�m�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�@���A����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��L���
�9�
�'�0�<����Y����V��C�U���%�b�0�l�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&ʹ��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��X�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ѓ�l_��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��
9��R	�����;�%�:�0�$�}�Z���YӖ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�8�N��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��R1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&Ĺ��
]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����֓�C9��S1�����&�<�;�%�8�8����T�����h��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�l�0�e�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ʹ��9��h��*���2�i�u�
���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�l�2�m����Y����T��E�����x�_�u�u���(߁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ӊ�
�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ց�&ù��l��G�����u�u�u�u�w�}�W���Y�����h��*���2�i�u�
���L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�l�0�f�<�(���&������^	�����0�&�u�x�w�}�����ד�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(ށ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����W����ߊu�u�u�u�w�}�W���Y���F��1��D���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�}�W���YӃ��Z �V�����1�
�e�|�#�8�W���Y���F�N��U���u�u�u�
���(�������A��S��*ӊ�
�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��L���d�%�0�u�$�4�Ϯ�����F�=N��U���
�
�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}�����ד�A��S��*ӊ�
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���R��Y��]���6�;�!�9�0�>�G������lV��h_�����l�
�%�1�9�t�^�����ƹF�N��U���u�u�9����4������� P��h��U��2�%�3�e�1�l�(���O�ԓ�C9��C��*��u�u�u�u�w�}�W�������W��R��!���0�=�&���.��������S��S�����
�
�
�e�1��N݁�	����F��UךU���u�u�u�u�w�}��������A��_��%���0��
�'������L���F��G1��E���d�
� �c�e�<�(�������l�N��U���u�u�u�3��2��������A��_��%���&�6�'�2�f�k�W������lV��h_�����l�
�%�'�#�/�(��Y���F�N��U����-��,�"��F�������F�	��*���b�c�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\���=�;�u�u�w�}�W���Y����_9��r*��6���!� �
�c�2�m����H����[��[1��0����:�!� ��k�G���I���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���`�3�8�d�~�<�ϰ��έ�l��D�����
�u�u�'���(���&����_��G1�����|�u�=�;�w�}�W���Y���F��[1�����0�8��&�6�8�4�������lW��E��D��u�h�2�%�1�m��������
9��h�� ���d�n�u�u�w�}�W���Y����_9��S������&�4�0��3����
����A��X�U��2�%�3�e�1�h����Mʹ��l��B��D��u�u�u�u�w�}�W�������W��R��6���4�0��;�%�1��������Q��S�����
�
�
�
�"�k�N���&����A��d��U���u�u�u�u�w�>�(�������^9��D�����;�'�9�&�e�/���N�����h��*���
� �c�l�6���������F�N��U���u�u�6�
�8�8����&����R��t�����&�f�'�2�f�e�W������lV��h[�� ��l�4�
�0�"�3�D�ԜY���F�N��Uʶ�
�:�0�!�%���������]��[1��A���2�d�m�u�j�:����I����l ��Z�����0� �;�a�]�}�W���Y���F�T�����!�'�
�4�4�9��������@9��E��D��u�h�2�%�1�m��������
9��h�� ���`�_�u�u�w�}�W���Y�Ư�l��R1�����4�6�1�1�8�)����&Ź��T9��V��Hʲ�%�3�e�3�b�;�(��&����V��Y1����u�u�u�u�w�}�W�������G��h-�����1�:�!�:���(���&����Z�P�����3�`�3�
�c���������]ǻN��U���u�u�u�u�;�3��������R��S�����:�
�
�
�2��A��E�ƫ�C9��1��@���
�a�
�%�%�)����B���F�N��U���u�9�;�1��8����
����W%��C��*���
�0�
�c�d�a�W���&����U9��Q��Aӊ�%�'�!�'��f�W���Y���F�N�����1�
�0�8��.����:����\
��h��*���m�i�u�'���(���&����_��G1�����
�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���˹��^9����U���}�4�
�:�$�����&���T��Q1�����3�
�e�
�'�9����P�Ƹ�VǻN��U���u�u�u�u��3��������Z��D=�����c�
�0�
�b�i�K�������9��1��*��
�%�'�!�%��L���Y���F�N��U���;�1�
�0�:�.����*����lW��h��*���e�i�u�'���(���&����_��G1�����
�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ޓ�@�� G��U���;�u�u�u�w�}�W���YӀ��K'��N!��*܊�0�
�c�`�k�}��������l��=N��U���u�u�u�u�w����� ����
9��P1�G���h�2�%�3��l�(��s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��ފ�&�
�|�|�#�8�}���Y���F�N�������g��#�o�(ށ�����Q�
N��*����g��!�e��(���H����CU��N��U���u�u�u�u�1��:���K����lT��1����d�u�h�3���;���6���� 9��Q��D���%�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9��G�����u�u�u�u�w�}�W�������f*��Y!��*���`�'�2�d�n�}�JϹ�	����T��G\�U���u�u�u�u�w�}����*����F��1�����d�e�u�h�0�-����Jǹ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�d�3�:�l�^�������F�N��U���u�u�3�
������&����Z��h_�����d�a�u�h�0�-����L˹��l�N��U���u�u�u�3���;�������_��[��*���
�`�c�i�w�/�(���N�ғ�]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��F���PӒ��]l�N��U���u�u�u�'�0�j�B��Y����U��X��G�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���܁�
����F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��D؊�&�
�d�|�~�)��ԜY���F�N��Uʧ�2�b�d�i�w�/�(���N�ԓ�]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����R��D��F���;�u�:�}�6�����&����P9��
N�����e�3�d�
�"�k�E���&����O�N���ߊu�u�u�u�w�}�W�������F�	��*���b�g�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y���R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����G^��D��\ʴ�1�;�!�}�'�>��������lV�	��*���
�
�
� �`�d�������F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��L���8�m�|�:�w�u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fځ�
����F��SN�����%�6�;�!�;�:���DӁ��l ��h��*���c�l�4�
�8�8�^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����_��D��M���|�!�0�_�w�}�W���Y���F��P1�@��u�'�
� �`�i���Y���F�N��U���0�
�l�u�j�:����&����CT��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�l�1�0�O������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���4�1�;�!��-��������Z��S�����
�
�
�
�"�k�N���&����O�N���ߊu�u�u�u�w�}�W�������F�	��*���b�a�%�n�w�}�W���Y���F��R	��E���h�2�%�3��h�(��s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���H����lW��G�����_�u�u�u�w�}�W���Y����W��S����� �b�a�%�l�}�W���Y���F���*��u�h�2�%�1��Cց�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϪ�ӈ��GF��V��]����
�&�|�8�}��������^��^ ��U���u�u�4�
��;����
����C��T�����&�u�4�
��;����	������h��*���e�3�
�l��-����UӁ��l ��h��*���b�l�4�
�8�8�W���&����U9��Q��Aӊ�%�1�;�y�6���������
OǻN�����_�u�u�u�w�<�Ͽ�&����@��Dd��U���u�u�u�"�2�}����&����U��N��U���u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����R��^	�����m�|�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���K����lW�	NךU���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y����[��V��!���f�3�8�g�j�}�W���Y���F�N�����
�&�u�h�6��#���M����lU��N��U���u�u�"�0�w�-�$���ǹ��^9��
P��U���u�u�u�u�w�}����*����Z�V��!���`�3�8�a�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N������3�8�i�w�-�$���Ź��^9��=N��U���u�u�u�=�9�<�(���
�Г�@��S����u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y�����YN��*���&�b�3�8�a�`�W���Y���F�N��U����
�&�u�j�<�(���
�ޓ�@��d��U���u�u�u�"�2�}����&����U�� N��U���u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y������T�����2�6�e�h�0�-�����ߓ�F9��1��*���0�|�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���@����l^�	NךU���u�u�u�u�w�}����&����[��G1��*���e�3�8�l�]�}�W���Y���D����&���!�e�3�8�n�`�W���Y���F�N��U����
�&�u�j�<�(���
����U��^�U���u�u�u�u� �8�W���*����W��D��E��u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d��.�(��s���F�N�����u�%��
�#�o����H���l�N��U���u�u�u�4������E�ƭ�l5��D�*���
�g�_�u�w�}�W���Y������d:�����3�8�d�u�i�W�W���Y���F�N��*���3�8�i�u�'��(���M����lW��=N��U���u�u�u�=�9�<�(���
����U��]��K�ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��h�����:�<�
�u�w�/�(���&����l ��W�����:�0�|�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����S��D��A�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��A���8�d�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GW��Q��D���k�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F��*���&�
�:�<��}�W���&����U9��Q��Aӊ�%�1�;�|�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�a�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��X�����`�h�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�<�(������F��h=����
�&�
�b�]�}�W���Y���D����&���!�m�3�8�f�}�I�ԜY���F�N��Uʴ�
��3�8�k�}����&����l ��h_����u�u�u�u�w�5�Ͽ�&����GW��Q��D���k�_�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�g�;���B���F�N��U���;�4�
��$�o�(���&���FǻN��U���u�u�u�u�'��(���Y����C9��h��D���8�g�n�u�w�}�W���Yӑ��]F��h=����
�&�
�e�j�}�W���Y���F�N�����
�&�u�h�6��#���K����^9��d��U���u�u�u�"�2�}����&����l ��h\�H���u�u�u�u�w�}�W�������l ��R������&�d�3�:�m�}���Y���F�@��U���0�&�h�u�]�}�W���Y���F�V��&���8�i�u����/���!����k>��o6��N���u�u�u�0�3�>���Y����]��E����_�u�u�x�6���������]F��X�����x�u�u�4��2����
����C��T�����&�}�%�6�{�<�(���&����l5��D�*���
�d�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�~�)����Y���F�N�����;�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����\��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��ʴ�&�2�u�'�4�.�Y��s���R��S�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������F�U�����u�u�u�<�w�u��������]��[����h�4�
�!�%�t�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\���=�;�_�u�w�}�W���Y����W
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��9���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������R��P �����&�{�x�_�w�}��������@��Y1�����u�'�6�&��-�������T9��R��!���g�
�&�
�f�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�o�^�������9F�N��U���u�%�'�4�.�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��m�DϿ�
����C��R��U���u�u�4�
�>�����I�Փ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��\�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�g�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���J�ƭ�@�������{�x�_�u�w�-��������U��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��D��u�h�}�%�4�3����H�����t=�����u�:�;�:�c�t�}���Y����C��R���ߊu�u�x�4��4�(���&������^	�����0�&�u�x�w�}��������W9��^�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����e�e�i�u�6�����&����F�V��&���8�d�u�:�9�2�F���B����������n�_�u�u�z�}��������lW��N�����u�'�6�&�y�p�}���Y����Z��S
��E���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�d�a�w�`�_�������l
��h_��U����
�&�}�n�9� ���Y���l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Cʴ�&�2�u�'�4�.�Y��s���R��^	�����e�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ފ�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����I���N��G1�����9�2�6�d�j�-�C���I����E
����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��[�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�����4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�F��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����T��V�����'�6�&�{�z�W�W���	����l��h_�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��o�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����0�g�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�d�d�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����M�ƭ�@�������{�x�_�u�w�-��������T��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ғ�lR��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�a�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1��A���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�F��Y����T��E�����x�_�u�u�'�.��������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�C���h�}�%�6�9�)����H����C9��h��]���:�;�:�d�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����L�ƭ�@�������{�x�_�u�w�-��������W��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ғ�lS��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�`�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1��@���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�F������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����d�e�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lR��hX�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��k�W�������A	��D�X�ߊu�u�%�&�0�?���@����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�C���N����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����V9��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�d�o�<����Y����V��C�U���4�
�<�
�3��@ׁ�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(߁�	����l�N�����u�u�u�u�w�}�W�������T9��S1�M��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�L����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�m�u�$�4�Ϯ�����F�=N��U���&�2�7�1�f�j��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�`�2�l������ƹF��R	�����u�u�u�u�w�}�W���
����W��Y��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ځ�&¹��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����d�c�4�&�0�}����
���l�N��*���
�1�
�l��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����_��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�h��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�g�`�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�`�0�f�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Aʴ�&�2�u�'�4�.�Y��s���R��^	�����d�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ߊ�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����H���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�`�0�c�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��]�����;�%�:�0�$�}�Z���YӇ��@��U
��G���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�����4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�E��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����U��V�����'�6�&�{�z�W�W���	����l��h\�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��n�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����0�c�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9�� 1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�g�f�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����L�ƭ�@�������{�x�_�u�w�-��������V��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ӓ�l^��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�`�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1��M���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����g�l�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lS��hW�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��k�W�������A	��D�X�ߊu�u�%�&�0�?���A����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�A���I����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����V9��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�`�<����Y����V��C�U���4�
�<�
�3��@؁�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(ށ�	����l�N�����u�u�u�u�w�}�W�������T9��S1�B��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�O����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�e�u�$�4�Ϯ�����F�=N��U���&�2�7�1�d�h��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�b�2�m������ƹF��R	�����u�u�u�u�w�}�W���
����W��[��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�&ù��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����f�a�4�&�0�}����
���l�N��*���
�1�
�d��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&���� W��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�f�f�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b�0�g�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Gʴ�&�2�u�'�4�.�Y��s���R��^	�����f�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*݊�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����J���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b�0�d�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��_�����;�%�:�0�$�}�Z���YӇ��@��U
��F���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�����4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�D��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&���� S��V�����'�6�&�{�z�W�W���	����l��h]�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��h�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����0�`�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�f�n�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����O�ƭ�@�������{�x�_�u�w�-��������^��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ѓ�lQ��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�c�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F�� 1��B���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�D������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����f�b�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lQ��hV�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��e�����Ƽ�\��D@��X���u�4�
�<��9�(�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������F�F��*���3�8�e�1� �)�W���DӇ��P	��C1��D��n�u�u�0�3�-����
��ƓF�C�����2�7�1�f�a�<����Y����V��C�U���4�
�<�
�3��Oف�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(ց�	����l�N�����u�u�u�u�w�}�W�������T9��S1�C��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�l�u�$�4�Ϯ�����F�=N��U���&�2�7�1�d�h��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�l�2�m������ƹF��R	�����u�u�u�u�w�}�W���
����W��[��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ց�&ù��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����a�a�4�&�0�}����
���l�N��*���
�1�
�e��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����V��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�a�f�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�d�
�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6��������� F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�f��(߁�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��A��4�&�2�u�%�>���T���F��h��*���
�f�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1�U���d�0�e�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
�f�8�G���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��A���&�<�;�%�8�8����T�����D�����a�e�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^���
�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�d���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Lʴ�&�2�u�'�4�.�Y��s���R��^	�����a�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*���0�g�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����M���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�d�2�o�������9F���U���6�&�n�_�w�}�Z���	����l��hZ�U���<�;�%�:�2�.�W��Y����C9��P1����m�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��Dۊ�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����L���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�d�
����������F�R �����0�&�_�_�w�}�ZϿ�&����Q��X����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����D���a�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���N�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�d�0�c�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W�� X�����;�%�:�0�$�}�Z���YӇ��@��U
��A���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�*���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�d�
�
��-����P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Mߊ�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��h_�����4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�C��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�d�0�c�6�����B����������n�_�u�u�z�}��������lR�������%�:�0�&�w�p�W�������T9��S1�C���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�a�c�i�w�<�(���
����9��
N��*���3�8�g�1� �)�W���B����������n�_�u�u�z�}��������lS�������%�:�0�&�w�p�W�������T9��S1�@���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�`�`�i�w�<�(���
����9��
N��*���3�8�c�1� �)�W���B����������n�_�u�u�z�}��������lS�������%�:�0�&�w�p�W�������T9��S1�A���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�`�a�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��Y�����;�%�:�0�$�}�Z���YӇ��@��U
��@���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�`�b�k�}��������_��N������3�8�d�w�2����H���9F���U���6�&�n�_�w�}�Z���	����l��h[�U���<�;�%�:�2�.�W��Y����C9��P1�����g�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�`�e�a�Wǿ�&����G9��1�Hʴ�
��3�8�`�9� ���Y���9F���U���6�&�n�_�w�}�Z���	����l��h[�U���<�;�%�:�2�.�W��Y����C9��P1�����a�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�`�c�a�Wǿ�&����G9��1�Hʴ�
��3�8�o�9� ���Y���9F���U���6�&�n�_�w�}�Z���	����l��h[�U���<�;�%�:�2�.�W��Y����C9��P1�����f�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�`�d�a�Wǿ�&����G9��1�Hʴ�
��3�8�f�}��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��B���&�<�;�%�8�8����T�����D�����`�c�4�&�0�����CӖ��P����6���&�|�u�u�5�:����Y���F�N��U���&�2�7�1�b�k�K�������]��[��D��4�
��3�:�l�W������O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�`�f�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�h�D��Yۇ��P	��C1��D��h�4�
��1�0�NϺ�����
O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�c�d�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�k�F��Yۇ��P	��C1��D��h�4�
��1�0�F�������W��UךU���;�u�'�6�$�f�}���Y���R��^	�����m�u�&�<�9�-����
���9F������7�1�c�l�6�.���������T��]���&�4�!�u���(߁�	����l��D��U���
�
�
�%�!�9��������lR��h\�����1�<�
�<�{�-�C���J����E
��^ �����%�a�0�a�6���������F��1��@���
�9�
�;�$�:�W���&����R��[
�����2�u�
�
����������@����*���
�%�#�1�>����	�ӓ�lW��G1�����
�<�y�%�b�8�E���&����Z��^	����0�f�4�
�;������Ƽ�9��1��*���
�;�&�2�w��(���&����_��Y1�����
�
�
�
�'�+����&������h��*���#�1�<�
�>�q�����ޓ�C9��S1��*���y�%�`�0�n�<�(���&����Z�G1�����4�
�9�
�9�.����&Ź��9��h��*���&�2�u�
���(�������]9��PB��*݊�
�
�%�#�3�4�(���UӖ��l��h�����<�
�<�y�'�j��������W9��h��Yʥ�b�0�a�4��1�(���
���C9��R1�����9�
�;�&�0�}�(؁�&Ź��l��h�����u�
�
�
��-��������TJ��hY��*Ҋ�%�#�1�<��4�[Ϯ�N����l��A�����<�y�%�l�2�m��������l��N��L���d�4�
�9��3����Y����l��h�����<�
�<�y�'�l�(���&����_��Y1�����
�d�0�d�6���������F��_��*؊�%�#�1�<��4�[Ϯ�H¹�� 9��h��*���&�2�u�
�f�8�C���&����Z��^	���
�
�
�%�!�9��������lW��R1�����9�
�;�&�0�W�W�������F�N��U���u�u�4�
�>�����A���N��h_�����4�
�9�
�9�.�������]��[����u�'�}�
�f�8�B���&����Z��^	��U���6�;�!�9�0�>�G����μ�W��hZ�����1�<�
�<�w�}��������\��h^�����%�d�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�H¹��9��h��*���&�2�h�4��2��������O��EN��*���0�d�4�
�;���������C9��Y�����6�e�u�'���F���I����E
��^ �����u�%�6�;�#�1����I�ƣ�N��^��*ڊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�l�2�l��������l��S�����;�!�9�2�4�m�W���Q����V9��V�����;�&�2�h�6�����&����P9����]���
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�@���A����E
��^ �����u�%�6�;�#�1����I�ƣ�N�� 1��B���
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
����������@��
N��*���&�
�:�<��t����	�ѓ�lS��G1�����
�<�u�u�'�>��������lV�X�����0�a�4�
�;���������C9��Y�����6�e�u�'���(���&����_��Y1����4�
�:�&��2����PӉ����h��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�b�0�f�<�(���&����Z������!�9�2�6�g�}����&Ĺ��9��h��*���&�2�h�4��2��������O��EN��*܊�
�
�%�#�3�4�(���Y�ƭ�l��D�����
�|�:�u�'�k��������W9��h��U���%�6�;�!�;�:���Y���C9��R1�����9�
�;�&�0�`��������_	��T1�U���}�
�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�L����l��A�����<�u�u�%�4�3��������F��F��@���c�4�
�9��3����DӇ��P	��C1�����e�u�'�}���(ځ�	����l��D��Hʴ�
�:�&�
�8�4�(�������lS��hZ�����1�<�
�<�w�}��������\��h^�����%�`�0�f�6���������[��G1�����9�2�6�e�w�/�_���&����R��[
�����2�h�4�
�8�.�(�������	����*���
�%�#�1�>�����Y����\��h�����|�:�u�%�b�8�G���&����Z��^	��U���6�;�!�9�0�>�G����μ�9�� 1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�
�'�+����&����F��h�����:�<�
�|�8�}�����ӓ�C9��S1��*���u�u�%�6�9�)�������\�G1�����4�
�9�
�9�.�������]��[����u�'�}�
���(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l��h�����<�
�<�u�w�-��������Z��N��U¥�a�0�d�4��1�(���
�����T�����2�6�e�u�%�u�(ہ�&ù��l��h�����h�4�
�:�$�����&����AF��G1�����h�4�
�:�$�����&���9F���U���6�&�n�_�w�}�Z���	����l��hY�U���<�;�%�:�2�.�W��Y����C9��P1����g�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�b�e�a�Wǿ�&����G9��1�Hʴ�
��3�8�d�9� ���Y���9F���U���6�&�n�_�w�}�Z���	����l��hV�U���<�;�%�:�2�.�W��Y����C9��P1����g�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�m�e�a�Wǿ�&����G9��1�Hʴ�
��3�8�f�}��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��D���&�<�;�%�8�8����T�����D�����l�d�4�&�0�����CӖ��P����6���&�|�u�u�5�:����Y���F�N��U���&�2�7�1�n�l�K�������]��[��D��4�
��3�:�l�W������O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h�����
�!�e�3�:�d�����Ƽ�\��D@��X���u�4�
�<��.����&����l ��hW�����;�%�:�u�w�/����Q����Z��S
��L���u�u�7�2�9�}�W���Yӏ����D�����`�f�u�=�9�W�W���Y���F��h��*���$��
�!�g�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	���&����
F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�d�1�0�F���
������T��[���_�u�u�%�$�:����&����GW��Q��Dڊ�&�<�;�%�8�}�W�������R��^	�����e�|�u�u�5�:����Y����������7�1�c�d�w�5��ԜY���F�N��*���
�&�$���)�F�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����l ��h_�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�E�������R��P �����&�{�x�_�w�}��������B9��h��G���8�d�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�d�~�}�Wϼ���ƹF�N�����%�&�2�7�3�h�C������F�N��U���4�
�<�
�$�,�$����ԓ�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��\�����d�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����Փ�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�f�3�8�f���������PF��G�����4�
�<�
�3��F���Y����V��=N��U���u�3�}�%�$�:����@���G��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�g�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*��4�&�2�u�%�>���T���F��h��*���$��
�!�c�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lS��N�����u�u�u�u�w�}��������V��c1��Dފ�&�
�f�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�d�
�$��D��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��Dߊ�&�
�a�4�$�:�W�������K��N�����<�
�&�$����������9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��C���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��i�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�d�
�&��h�����Ƽ�\��D@��X���u�4�
�<��.����&����l ��h_�����2�
�'�6�m�-����
ۇ��@��U
��D��|�u�u�7�0�3�W���Y����UF��G1�����1�d�a�|�#�8�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
����U��[��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�l�(���&����@��YN�����&�u�x�u�w�<�(���&����l5��D�*���
�b�4�&�0�����CӖ��P�������7�1�m�g�]�}�W������F�N��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���%�&�2�6�2��#���H˹��^9��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���Hʹ��^9�������%�:�0�&�w�p�W�������T9��R��!���d�
�&�
�o�<����&����\��E�����%�&�2�7�3�h�A�ԜY�Ʈ�T��N��U���<�u�4�
�>�����N����[��=N��U���u�u�u�%�$�:����&����GW��Q��D���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GW��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�d�3�:�m��������\������}�%�&�2�5�9�D���Y����V��=N��U���u�3�}�%�$�:����J����[��=N��U���u�u�u�%�$�:����&����GW��D��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��W�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�g�
�&��d��������\������}�%�&�2�5�9�F��P�����^ ךU���u�u�3�}�'�.��������O��_�����u�u�u�u�w�-��������`2��C\�����d�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�e�3�8�f�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C\�����g�u�&�<�9�-����
���9F������6�0�
��$�o�(���&�ד�@��Y1�����u�'�6�&��-��������T��=N��U���<�_�u�u�w�}����	����l��h_�F���=�;�_�u�w�}�W���Y����Z��D��&���!�g�3�8�e�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�o����K�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���K����lW��D�����:�u�u�'�4�.�_���
����W��X����u�0�<�_�w�}�W����έ�l��h��*��b�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���J����lT��D�����:�u�u�'�4�.�_���
����W��X��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��A��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lQ��d��Uʷ�2�;�u�u�w�}��������T9��S1�G���=�;�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ߊ�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�B����ғ�@��Y1�����u�'�6�&��-��������U��=N��U���<�_�u�u�w�}����	����l��h_�F���=�;�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��݊�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�@����Г�@��Y1�����u�'�6�&��-��������S�N�����;�u�u�u�w�4�Wǿ�&����Q��^�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��*���
�u�&�<�9�-����
���9F������6�0�
��$�e����N����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:��Ҋ�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��CW�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�n�;��������]9��X��U���6�&�}�%�$�:����L���F�U�����u�u�u�<�w�<�(���&����S�����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u��-��$����N�ד�F9��[��D��u��-� ��3����J�ӓ�V��W����u��-��.�(�(�������9��R�����b�`�_�u�w�����-����G9��h_�� ��e�
�f�i�w�}�W���YӀ��K+��c\�� ���f�3�
�m��l� ���Yە��l��1�����e�d�%�}�~�`�P���Y����l�N��Uʧ�2�b�`�_�w�}�$���,����|��]��*���d�b�
�d�k�}�(�������9��h_�G���n�u�u�3���;���6���� 9��Q��D���%�u�h�_�w�}�W���*����2��x��Gي�
� �d�b��l� ���Yە��l��1��*���d�l�
�g�g�}�W��PӃ��VFǻN��U����-� ��9�(�(���L����lW��UךU����-� ��9�(�(�������9��R�����&�9�
�a�1��@܁�L���F��h��9����!�g�
�9�8����H����
W��G\��Hʦ�1�9�2�6�!�>����������T�����d�
���~�v�����μ�a��[��*���l�`�%�|�l�}�Wϸ�&����gT��B��F���
�-�
�
��(�F��&���F��S1�����#�6�:�}�>�3�ǿ�&����G9��V��3���|�~�&�2�2�u�(�������9��h_�A���|�n�u�u�1��:���K����lT��^ �����0�d�3�
�g�k����D���F�N�����<�<�<�e�4�.�(�������V��h����u�&�9�!�'��D���&����l��G��U��|�0�&�u�w�}�W���
����^��1��*��c�%�n�u�w�;�(���5�Ԣ�F��1��*���,�0�3�
�n��D��Y���F���*؊�
�
�
�4�#�>��������l��@��U¦�9�!�%�
��(�O���	����[�I�����u�u�u�u�w�.����	����F9�� 1��N�ߊu�u�x�2�'�;�G���Hù��lP��h�����&�<�;�%�8�8����T�����h��*���e�3�
�l��-����
����l��TN����0�&�4�
�2�}��������B9��h��A���8�d�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�u�'��-��������Z��S�����2�6�0�
��.�F܁�
����O����ߊu�u�u�u�w�}����&ù��V��B1�G���
�0�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӁ��l ��h��E���
�l�
�%�4�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�'���(���I����_��V�����u�h�2�%�1�m���&����
T��G1�����4�
�!�'��8�L���YӁ��l ��h��E���
�l�
�;��4�2�������A��[��Hʥ�c�0�e�<��4�L���YӁ��l ��h��E���
�l�
�;������&˹��F���*���
�;�&�2�]�}�W���&����U9��h��C���<�
��2�>�.�O���H���C9��R1�����<�n�u�u�0�-��������U��\������4�2�
���W��	�ӓ�lV��Y1���ߊu�u�'�
���(�������9��h>�����0�l�0�d�k�}�(ځ�&¹��l��d��Uʲ�%�3�e�3�f����K����`��R'��E���e�i�u�9���5�������G9��h��*���
�`�b�_�w�}����&ù��V��B1�G���
�$�f�i�w�8�(��B�����h��*���e�3�
�l��3����Y����lP��h_�����2�_�u�u�%��(߁�&�֓�F9��1��*���0�
�u�h�'�d��������T]ǑN��X���'�
�
�
�����@����P��D��ʥ�:�0�&�u�z�}�WϹ�	����l ��h��C���4�
�0�4�$�:�(�������A	��D�����y�4�
�<��.����&����l ��h_�U���
�
�
�
�g�;�(��&����\�������6�0�
��$�l�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�u��������_	��T1�Hʴ�
�<�
�&�&��(���M����lW����U���}�4�
�:�$�����&���T��Q1����
� �c�g�6�����P�ƣ�N��h�����:�<�
�u�w�-��������`2��C_�����d�|�|�u�?�3�}���Y���F�P�����3�`�3�
�c�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʲ�%�3�e�3�b�;�(��&����VF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����U9��Q1�����a�
�%�&�6�)�K�������9��1��*��
�%�&�4�#�<�(�������T]ǻN�����
�
�
�
�"�k�N���&����@9��R1�I���
�
�
�
�9�.��ԜY�ƫ�C9��1��@���
�a�
�;��4�������F�� 1��F���
�<�n�u�w�:����I����l ��Z�����4�;�
�
��}�JϮ�N����l��D�����u�'�
�
���(���O�ߓ�]9��^ ��A���f�i�u�
���(���
����F�P�����3�`�3�
�c���������l��R�����0�c�<�
�>�f�W�������lV��h[�� ��l�<�
�4�9��(���Y����lQ��hY�����2�_�u�u�%��(߁�&ƹ��lP��h��2���&�a�0�c�k�}�(؁�&˹��l��d��Uʲ�%�3�e�3�b�;�(��&����R��hZ��*���h�%�b�0�n�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�g�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�f�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�e�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�d�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�c�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�b�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�a�4�(���B�����h��*���
� �c�l�>���������A	��\��*���h�%�a�0�`�4�(���B�����h��*���
� �c�l�>��!������F��h �����'�
�=�0��<����&����A��[�N���u�2�%�3�g�;�B���&����Z��a1����i�u�
�d�2�k������ƹF��E��*ڊ�
�
� �c�n�4�(���K����Z�Q=��4����!�g�
�2��B��s���T��Q1�����3�
�a�
�9��(݁�&�����hY�N���u�2�%�3�g�;�B���&����Z��V ��*݊�
�u�h�%�b�8�E���&����9F�	��*���
�
�
� �a�d��������9��N�U���
�
�
�;�$�:�}���Y����U9��Q1�����a�
�;��9�8�@���K���C9��R1�����<�n�u�u�0�-�����ӓ�F9��1��*���2�
�
�
�w�`�����ӓ�]9��PUךU���'�
�
�
�����@����a��R1����i�u�
�
���������F��G1��E���`�3�
�a��3�%����ѓ�lS�
N��@���b�<�
�<�l�}�WϹ�	����l ��h��C���<�
�4�2���(���DӖ��l��h�����_�u�u�'���(���&����_��Y1�����b�0�b�i�w��(���&����Z��N�����3�e�3�`�1��Cց�����9��N�U���
�
�
�;�$�:�}���Y����U9��Q1�����a�
�;����(���DӖ��9��1��*���n�u�u�2�'�;�G���L����R��^ �����
�u�h�%�n�8�F���&����9l�N�U���
�
�
�
��(�@���������^	�����0�&�u�x�w�}�����֓�l_��B1�L���
�0�4�&�0�����CӖ��P�������4�
�<�
�$�,�$���Ĺ��^9�������6�0�
��$�e����N���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u��-��������Z��S�����2�6�0�
��.�@������\�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�u�?�3�}���Y���F�P�����3�l�3�
�g�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʲ�%�3�e�3�n�;�(��&����VF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����U9��Q1�����e�
�%�&�6�)�K�������9��1��*��
�%�&�4�#�<�(�������T]ǻN�����
�
�
�
�"�j�N���&����[��[1��0����:�!� ��k��������W��=d��U���u�'�
� �`�k����
������T��[���_�u�u�'��(�@�������@��h����%�:�0�&�6�����
����g9��1����u�%�6�y�6�����
����g9��Z�����f�u�'�
���(�������9��h
�����%�&�2�6�2��#���A����lQ�V�����&�$��
�#�����UӇ��@��T��*���&�d�
�&��i�W���
����@��d:�����3�8�d�y�6���������
J��G1�����0�
��&�c�;���s���Q��Yd��U���u�<�u�}�8�u��������_	��T1�Hʴ�
�0�|�:�w�<�(���
����T��N�����<�
�&�$���ׁ�
����	�������!�9�2�6�f�`��������V��c1��L���8�m�u�'��-��������Z��S�����2�6�0�
��.�Fځ�
����F��F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�8�}��������_	��T1�Hʴ�
�<�
�&�&��(���&���� O��EN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9��������W9��G�����4�
�:�&��2����Y�ƭ�l��h�����
�!�a�3�:�l�^Ͽ��έ�l��D�����
�u�u�'���(���I����_��V�����|�|�!�0�w�}�W���Y�����h��B���6�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����U��X����u�%�6�;�#�1����H���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����3�
�d�
�'�2�Ͽ�
����C��R��U���u�u�2�%�1��Fف�	����l��^	�����u�u�'�6�$�u��������B9��h��*���
�y�4�
�>�����*����T��D��D���%�&�2�6�2��#���Hù��^9�������7�1�c�l�w�-��������`2��C[�����y�4�
�<��.����&����l ��h_�U���&�2�6�0��	���&����_�N�����;�u�u�u�w�4�W�������]��[����h�4�
�<��.����&����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��h�^������F�N��U���2�%�3�
�f��������R��X ��*���
�n�u�u�w�}�������R��X ��*���<�
�u�u�'�.��������l��1����|�:�u�4��2��������F�V�����&�$��
�#�m����@�ƣ�N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�8�u��������lP��G�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��d�^������F�N��U���2�%�3�
�f��������R��X ��*���
�n�u�u�w�}����Y���F�N��U���
� �b�c�8�>����D�Ĕ�]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�'�
� �`�k����
������T��[���_�u�u�'��(�@���	ù��@��h����%�:�0�&�6�����
����g9��1����u�
�d�0�d�4�(���UӖ��9��1��*���y�4�
�<��.����&����l ��h_�U���
�l�y�'�0�e�F���	����l��F1��*���e�3�8�l�w�����-����l+��C�����'�2�d�f�{�<�(���&����l5��D�����a�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���I����lW��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������F9��1��U��'�2�b�f�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��G���8�d�|�u�?�3�}���Y���F�P�����d�
�e�i�w�����-����l+��C�����'�2�d�f�l�}�W���YӃ��Z �F��*���&�
�:�<��}�W���
����@��d:�����3�8�l�u�%�u��������\��h_��U���&�2�6�0��	���&����S�N�����u�u�u�u�w�}��������9��R�����m�d�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y�ƫ�C9��hY�*��i�u�
�d�2�n������ƹF�N�����u�}�%�6�9�)���������D�����
��&�d�1�0�G�������9F�N��U���u�'�
� �`�k����DӖ��9��1��*���n�u�u�u�w�8����Y���F�N����� �b�c�%�w�`�U���!����k>��o6��-���������U�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�P�����d�
�d�4�$�:�W�������K��N�����3�
�d�
�f�<����&����\��E�����%�&�2�6�2��#���H����lV�G1�*���
�;�&�2�w�-��������`2��C_�����d�y�'�2�`�h�W���&������D�����
��&�d��.�(������f*��Y!��*���d�'�2�d�g�q��������V��c1��@���8�a�u�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����֓�@��GךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���!�0�u�u�w�}�W���YӁ��l �� _�����h�'�2�m�f�W�W���Y�Ʃ�@��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�|�8�}��������_	��T1�Hʴ�
�<�
�&�&��(���O����lW����]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�n�t�W������F�N��Uʲ�%�3�
�d��l�K�������]ǻN��U���9�<�u�}�'�>��������lW������6�0�
��$�h����M����[��=N��U���u�u�u�'��(�@���	��� ��O#��!ػ� �
�f�d�%�:�F��B���F������}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�^Ϫ���ƹF�N��U���'�
� �b�a�-�W��	����V9��^ ����u�u�u�u�2�.�W���Y���F�	��*���b�c�%�u�j��/���!����k>��o6��-���������}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��G1��*��
�0�4�&�0�}����
���l�N�����
�g�
�0�6�.���������T��]���&�2�6�0��	��������F��h��U���&�2�6�0��	���&����U�P�����3�d�
� �a�o�������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�m�u�'�.��������l��1����y�4�
�<��.����&����l ��h_�U���&�2�7�1�a�d�W���
����@��d:��ފ�&�
�|�u�w�?����Y���F��QN�����}�%�6�;�#�1����H����C9��G�����%�6�;�!�;�:���DӇ��@��T��*���&�m�3�8�`�}����	����@��X	��*���u�%�&�2�4�8�(���
�ߓ�@��N��U´�
�:�&�
�8�4�(���Y����Z��D��&���!�`�3�8�f�t��������]��[����h�4�
�<��.����&����l ��h_�U���}�%�6�;�#�1����H����C9��P1������&�a�3�:�n�W���Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�%�&�2�5�9�A��Y�����T�����2�6�d�h�6�����
����g9��Z�����f�u�;�u�6�����&����P9��
N�����e�3�d�
�"�k�E���&����O����ߊu�u�u�u�w�}��������l��S�����;�!�9�2�4�m�}���Y���V
��d��U���u�u�u�2�'�;�(��&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӁ��l �� \�����1�u�&�<�9�-����
���9F�	��*���b�g�:�6�3���������PF��G�����4�
�<�
�$�,�$���¹��^9�������6�0�
��$�l�(���&���R��^	������
�!�e�1�0�N���	����l��hX�Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�f�����L�ƭ�l��h�����
�!�e�3�:�l�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1�����0�
��&�f�����H�ƣ�N��h�����:�<�
�u�w�-��������`2��C_�����l�u�'�}�6�����&����P9��
N��*���
�&�$���)�(���&����]��X�����2�7�1�c�n�t��������]��[����h�4�
�<��.����&����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��d�^������F�N��U���2�%�3�
�e��������R��X ��*���
�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��h��*���|�!�0�u�w�}�W���Y����A��B1�G���6�1�u�h�6�����&����]ǻN��U���9�0�_�u�w�}�W���Y����U��\�����0�i�u��u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���T��Q��G؊�e�4�&�2�w�/����W���F�P�����g�
�e�4�$�:�(�������A	��D�����2�6�0�
��.�F������C9��h��*���&�2�u�
�f�8�C���&������D�����
��&�d��.�(��Y����_�������6�0�
��$�l�(���&����V��V����<�
�&�$���ځ�
������D�����
��&�d��.�(��Y����Z��D��&���!�e�3�8�f�t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�g�1�0�F���Y����l�N��U���u�2�%�3��o�(��E�ƾ�T9��UךU���u�u�9�<�w�u��������_	��T1�Hʴ�
�<�
�&�&��(���I����l_�X�����:�&�
�:�>��W���	����l��F1��*���c�3�8�d�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����֓�@��G��U���;�_�u�u�w�}�W�������lQ��h�I���0�
�l�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�����a�|�!�0�w�}�W���Y�����h��B���%�u�h�%�f��(߁�����l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�2�%�1��E݁�I���C9��h��*���&�2�_�u�w�}�W������F�N��Uʲ�%�3�
�g��m�K���!����k>��o6��-���������/���B���F���U���u�u�u�0�3�-����
��ƓF�C����� �b�g�%�w�.����	����@�CךU���'�
� �b�e�-�(�������A	��N�����&�4�
�<��.����&����U��B��*���0�`�<�
�>�q��������V��c1��D؊�&�
�d�u�2��O������P�V�����&�$��
�#�m����@�ƪ�l��{:��:���g�
�
�0��h�E���*����2��B�� ���%�,�d�
�2��B��Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�*���
�`�u�%�$�:����&����GT��Q��D���u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C\�����d�|�u�=�9�W�W���Y���F��G1��*��
�d�i�u�2��O��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��l�^Ϫ���ƹF�N��U���'�
� �b�e�-�W������f*��x��8���<�9�
�`�%�:�F��B���F������}�4�
�:�$�����&���R��^	������
�!�e�1�0�N����έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�!�0�u�w�}�W���Y����A��B1�G���u�h�'�2�o�k�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����
�g�
�d�k�}�$���,����|��]��*���
�`�g�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C_�����|�u�=�;�]�}�W���Y���T��Q��G؊�d�i�u�
�f�8�B���&����9F�N��U���0�_�u�u�w�}�W�������lQ��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������9�������%�:�0�&�w�p�W�������F9��1��*���<�;�%�:�w�}����
�έ�l��h�����
�!�
�&��q�����ƭ�l��h�����
�!�
�&��q��������W9��B�����2�6�0�
��.�E������F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�u��������\��h_��U���&�2�6�0��	��������F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}����	����l��hX�\���'�}�%�6�9�)���������D�����
��&�g�1�0�F���PӒ��]FǻN��U���u�u�'�
�"�j�O���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʲ�%�3�
�g��8�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�:����&����P��D��ʥ�:�0�&�u�z�}�WϹ�	����U��T�����;�%�:�u�w�/����Q����Z��D��&���!�
�&�
�{�<�(���Y����Z��D��&���!�
�&�
�{�<�(���&����^�������6�0�
��$�o����H���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u��-��������Z��S�����2�6�0�
��.�D������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�2�_���
����W��W��U���}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�^�������9F�N��U���u�'�
� �`�i����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����3�
�f�
�2�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�0�-����Mǹ����^	�����0�&�u�x�w�}��������9��h�����%�:�u�u�%�>��������J��R	��M���4�
�<�
�$�,�$���˹��^9�������6�0�
��$�d����A�ƭ�l��h�����
�!�`�3�:�l�[Ͽ�&����P��h=����
�&�
�m�w�8�(��UӇ��@��T��*���&�d�
�&��q��������V��c1��Dۊ�&�
�e�u��%�"�������lT��R	��@��u��-� �.�(�(ց�����^�Q=��4����!�c�'�0�l�D������lV��h[�� ��l�4�
�0�"�3�F������T9��R��!���g�
�&�
�f�W�W�������F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��F�������9F�N��U���u�'�
� �`�i����DӀ��K5��N!��*ӊ�0�
�c�m�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��L���8�d�|�u�?�3�}���Y���F�P�����a�
�e�i�w����� ����9��P1�F��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������F9��1��U��2�%�3�e�1�h����Mʹ��l��B��D��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������F9��1��U��'�2�m�d�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��E���8�l�|�!�2�}�W���Y���F��E�� ��a�%�u�h�%�:�@��s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��Uʲ�%�3�
�a��m�K�������]ǻN��U���9�<�u�}�'�>��������lW������6�0�
��$�e����N����[��=N��U���u�u�u�'��(�@���	��� ��O=�����
�e�g�'�0�l�G��Y���F��[�����u�u�u�u�w�/�(���N�ғ�F�L��-���������/���!����k>��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�2�'�;�(��&����@��YN�����&�u�x�u�w�:����&����CW��D�����:�u�u�'�4�.�_���
����@��d:��Ҋ�&�
�y�4��4�(�������@��Q��M���%�&�2�6�2��#���Hƹ��^9��N��*���
�&�$���)�N���������D�����
��&�d��.�(������T9��R��!���d�
�&�
�g�}�$�������A��^ �����#�
�c�
�2��B��Y����Z��D��&���!�g�3�8�e�t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�g�1�0�E���Y����l�N��U���u�2�%�3��i�(��E�ƭ�l��D�����f�`�e��l�}�W���YӃ��Z �F��*���&�
�:�<��}�W���
����@��d:��ӊ�&�
�|�:�w�<�(���
����T��N�����<�
�&�$����������O��EN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�e�~�}����s���F�N�����3�
�a�
�f�a�W�������G��h������#�
�c��8�(��M���F�N�����}�}�%�6�9�)���������D�����
��&�m�1�0�@����έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���:�u�4�
�8�.�(�������F��h��*���$��
�!�g�;���P�Ƹ�V�N��U���u�u�2�%�1��Cہ�H���R��X ��*���g�f�f�e��f�W���Y����_��=N��U���u�u�u�'��(�@���	���D��o6��-���������/���!����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�2�%�3��i�(������]F��X�����x�u�u�2�'�;�(��&�֓�@��Y1�����u�'�6�&��8�(��UӔ��lQ��N����`�u�%�&�0�>����-����l ��hY����<�
�&�$���ց�
������D�����
��&�d��.�(��Y����Z��D��&���!�l�3�8�f�q����A���R��^	������
�!�e�1�0�N���	����l��F1��*���d�3�8�d�{�;�(���;����l_��R	��C��u�'�
�
���(���O�ߓ�C9��C��*��_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�m�|�!�2�}�W���Y���F��E�� ��l�%�u�h�1��$���6����l��h_�M�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��Z��U���;�_�u�u�w�}�W�������lQ��h�I���'�
�
�
�����@����A��E ��D�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��^��U���;�_�u�u�w�}�W�������lQ��h�I���0�
�d�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�|�u�=�9�W�W���Y���F��G1��*��
�e�i�u�2��A��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�l�3�8�o�t����Y���F�N��U���
� �b�l�'�}�JϬ�����l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�2�%�1��Cց�I���A�� Y����u�u�u�9�2�W�W���Y���F��G1��*��
�e�i�u���/���!����k>��o6��-�������l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����A��B1�L���u�&�<�;�'�2����Y��ƹF��E�� ��l�%�
�&�>�3����Y�Ƽ�\��DF��*���
�&�$���)�(���&����C9��P1������&�l�3�:�e�W���
����@��d:�����3�8�d�y�6�����
����g9��W�����m�u�%�&�0�>����-����9��Z1�U���&�2�6�0��	���&����V�Q=�����!�'�
�<�4�.�0���&����A��[�\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���T��Q��Aӊ�d�i�u�%�4�3����J����wW��r\�U���u�u�0�&�1�u�_�������l
��^��U���%�&�2�6�2��#���@����l^�X�����:�&�
�:�>��W���	����l��F1��*���`�3�8�d�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ד�@��G��U���;�_�u�u�w�}�W�������lQ��h�I����;�1�
�2�0��������E��V�����`�e�_�u�w�}�W��������T�����2�6�d�h�6�����
����g9��1����u�'�}�%�4�3��������[��G1�����0�
��&�f�����P����[��=N��U���u�u�u�'��(�@���	�����T�����f�
��d�b�n�}���Y���V
��d��U���u�u�u�2�'�;�(��&���F��o6��-���������/���!����k>�=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�'�
�"�j�C���Y����T��E�����x�_�u�u�%����M����R��P �����o�%�:�0�$�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1�Yʧ�2�b�f�u�'�.��������l��1����y�'�2�m�o�}����&ù��9��hX�*���'�!�'�
�g�W�W�������F�N�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��C�������9F�N��U���u�'�
� �`�i����DӁ��l ��h��*���c�l�4�
�2�(���B���F������}�%�6�;�#�1����H����C9��P1������&�d�
�$��G�������9F�N��U���u�'�
� �`�i����DӔ��l^��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���ց�
����F��R ��U���u�u�u�u�0�-����Lǹ��Z�E��B��_�u�u�u�w�1��ԜY���F�N�����
�`�
�e�k�}�/���!����k>��o6��-���������L���Y�������U���u�0�1�%�8�8��Զs���K��E�� ��m�%�u�&�>�3�������KǻN����� �b�m�%��.����	����	F��X��´�
�<�
�&�&��(���&����J��G1�����0�
��&�f�����M�ƾ�T9��B�����2�6�0�
��.�Fށ�
����F��P1�M���'�
�
�
�����@����A��E ��E�ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�6�����
����g9��[�����a�|�!�0�w�}�W���Y�����h��B���%�u�h�2�'�;�G���L����R��V�����;�d�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��_�����e�|�!�0�w�}�W���Y�����h��B���%�u�h�'�0�e�O�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����3�
�`�
�g�a�W���&����9F�N��U���0�_�u�u�w�}�W�������lQ��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�;�>�!��&���� _��N�U���-��,� ��j����Kƹ��T��N����!�u�|�_�w�}����&�֓�F9��V��A��u��-��.�(�(���H����V��h�F���:�;�:�g�~�W�W�������W��B1�GҊ�d�i�u��/�����&�ѓ�l ��^�*��g�u�u�u�8�3���B���
��h8�� ��l�%�u�h�1��6���6����9��hV�*��f�u�:�;�8�o�^�ԜY�Ƽ�T��h_��D���
�d�c�%�w�`�}���Y���R��X ��*���f�e�"�0�w�)���&����T��G\��\��r�r�u�9�2�W�W���Y�Ơ�P9��_�� ��g�
�d�_�w�}�(��I�ד�l ��]�����h�_�u�u�w�}��������ET��N�����!�%�&�3��n�(��I���W����ߊu�u�u�u�8��(�������
9��d��Uʥ�e�0�e�i�w�1����&����l2��R������
�'�
��8�(��K��ƹF�N��E���e�4�
�9�w�.����	����@�CךU���
�
�
�
�'�+����
����C��T�����&�}�%�6�{�<�(���&����l5��D�*���
�d�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�g�|�~�)����Y���F�N��*ڊ�
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��h^��*ڊ�%�#�1�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%�e�0�d�k�}��������A��_��%���0��
�'������L����9F�C����0�d�4�
�;�}����Ӗ��P��N����u�
�
�
��-��������]9��X��U���6�&�}�%�4�q��������V��c1��G؊�&�
�d�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���g�3�8�g�~�t����Y���F�N��U���
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���*���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�e�0�e�a�W�������G��h-�����1�:�!�:������L����9F�C����0�g�4�
�;�}����Ӗ��P��N����u�
�
�
��-��������]9��X��U���6�&�}�%�4�q��������V��c1��G؊�&�
�d�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���g�3�8�g�~�t����Y���F�N��U���
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���*���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�e�0�d�a�W�������G��h-�����1�:�!�:���(���&����lǻN��Xʥ�e�0�f�4��1�W�������A	��D�X�ߊu�u�
�
����������Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�d�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�e�t�^Ϫ���ƹF�N��U���
�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8����Y���F�N��*ڊ�
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�e�2�i�K�������V9��E�����1�1�:�!�8��(݁�����^��=N��U���%�e�0�a�6�����
������T��[���_�u�u�
���(�������@��Y1�����u�'�6�&��-�������T9��R��!���g�
�&�
�f�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�o�^�������9F�N��U���u�
�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�%�g�8�B��Y����\��C��*���6�1�1�:�#�2�(���&����S��dךU���x�%�e�0�b�<�(���Y����T��E�����x�_�u�u���(ځ�	����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�g�
�&��l�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�g�1�0�E���PӒ��]FǻN��U���u�u�
�
���������R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�m���E�Ư�l��R1�����4�6�1�1�8�)����&ǹ��T9��V����u�x�%�e�2�k�����ƭ�@�������{�x�_�u�w��(���&����_��D�����:�u�u�'�4�.�_�������C9��P1������&�g�
�$��F�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�e�;���P����[��=N��U���u�u�u�
���(������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�
�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�-�G���N���P
��X
�����
�4�6�1�3�2����&����A��[�N�ߊu�u�x�%�g�8�@���&����R��P �����&�{�x�_�w�}�(߁�&Ĺ��l��h�����%�:�u�u�%�>����	������D�����
��&�g��.�(��s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�o����K�����YNךU���u�u�u�u���(؁�	����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�
���������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}�������F��h �����'�
�4�6�3�9��������9��P1�L��_�u�u�x�'�m��������WF��D��U���6�&�{�x�]�}�W���&����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�����H���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�E�������O��_�����u�u�u�u�w��(���&����_�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�
���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�I����Z�T�����!�'�
�4�4�9��������@9��E��D��n�_�u�u�z�-�G���@����E
��V�����'�6�&�{�z�W�W���&ù��
9��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�o�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O����ߊu�u�u�u�w�}�(߁�&ʹ��l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u���(ց�	����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lW��R1�����9�
�;�&�0�<����Y����V��C�U���%�d�
�
��-��������T9��D��*���6�o�%�:�2�.���&����R��[
���
�
�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��Dڊ�
�
�%�#�3�t����Y���F�N��U���e�0�e�4��1�(���
���F��^��*ڊ�%�#�1�_�w�}�W������F�N��U���%�d�
�
��-��������TF���E���e�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�*���
�;�&�2�6�.��������@H�d��Uʥ�d�
�
�
�9�.����
����C��T�����&�}�
�e�2�m�W���I����l��PB��*���0�e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��h��*���#�1�|�!�2�}�W���Y���F��h_�����<�
�<�u�j�-�F߁�&��ƹF�N�����_�u�u�u�w�}�W���I����l��D��I���
�e�0�e�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h_�����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�d���(�������]9��P1�����
�'�6�o�'�2����	����V9��V�����%�d�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�d�
�
�
�'�+��������9F�N��U���u�
�d�0�g�<�(���&����Z�
N��Dۊ�
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�d���(�������]9��PN�U���d�0�e�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�d�
����������Z��G��U���'�6�&�}��l���Y����l��h�����
�d�0�e�6�����Y����V��=N��U���u�3�}�4��2��������F�G1�*���
�%�#�1�~�)����Y���F�N��*���0�e�<�
�>�}�JϮ�H¹��]ǻN��U���9�0�_�u�w�}�W���Y����l��h�����i�u�
�d�2�m����B���F���U���u�u�u�0�3�-����
��ƓF�C��*���0�d�4�
�;�����Ӈ��Z��G�����u�x�u�u�'�l�(���&����_��Y1�����&�2�
�'�4�g��������lW��R1�����9�y�%�d���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�d�
����������[��=N��U���u�u�u�
�f�8�F���&����Z��^	��Hʥ�d�
�
�
�'�+��ԜY���F��D��U���u�u�u�u�'�l�(���&����_��Y1����u�
�d�0�f�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�d�
�
��3��������]F��X�����x�u�u�%�f��(ށ�����l��^	�����u�u�'�6�$�u�(������C9��h��*���2�u�
�d�2�l������ƹF��R	�����u�u�u�3��<�(���
����T��N����
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�d�0�d�>�����DӖ��9��UךU���u�u�9�0�]�}�W���Y���C9��h��*���&�2�i�u��l����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�d�0�g�6�����������^	�����0�&�u�x�w�}���&����R��[
�����2�4�&�2��/���	����@��h_�����4�
�9�y�'�l�(���&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�f��(݁�	����O��_�����u�u�u�u�w��F���K����E
��^ �����h�%�d�
���������F�N�����u�u�u�u�w�}���&����R��[
�����2�i�u�
�f�8�E���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�d���(���
����@��YN�����&�u�x�u�w�-�Fށ�&����l��h�����%�:�u�u�%�>����&�ד�lT�G1�*���
�'�2�u��l��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�d�
�
��-����PӒ��]FǻN��U���u�u�
�d�2�o���������1��G�ߊu�u�u�u�;�8�}���Y���F�G1�*���
�;�&�2�k�}�(����ԓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�d�2�n��������l�������%�:�0�&�w�p�W���	����V9��V�����;�&�2�4�$�:�(�������A	��D��*���0�f�4�
�;�q���&����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�Fށ�&����l��G�����_�u�u�u�w�}�W���H����l��A�����<�u�h�%�f��(܁�	����l�N��Uʰ�&�u�u�u�w�}�W���	����V9��V�����;�&�2�i�w��F���J����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�l�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�H¹�� 9��h��*���<�;�%�:�w�}����
�μ�W��h]���
�
�
�'�0�}�(����Փ�C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�d���(��������YNךU���u�u�u�u��l��������TF���D���f�_�u�u�w�}����s���F�N����
�
�
�;�$�:�K���&�ד�lU��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u��l��������W9��h��U���<�;�%�:�2�.�W��Y����lW��R1�����9�
�;�&�0�<����&����\��E�����
�d�0�a�6����	����V9��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�H¹��9��h��\���=�;�_�u�w�}�W���Y����l��h�����<�
�<�u�j�-�Fށ�&ǹ��l��d��U���u�0�&�u�w�}�W���Y����lW��R1�����9�
�;�&�0�a�W���H����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��9��1��*���
�&�<�;�'�2�W�������@N��_��*���%�d�
�
��/����&�ד�lR��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�l�(���&����_����ߊu�u�u�u�w�}�(����ғ�]9��PN�U���d�0�a�_�w�}�W������F�N��U���%�d�
�
��3����E�Ƽ�W��hZ�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(����ӓ�C9��S1��*���u�&�<�;�'�2����Y��ƹF��h_�����4�
�9�
�9�.����
����C��T�����&�}�
�d�2�h��������lW��R1�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��9��1��*���|�u�=�;�]�}�W���Y���C9��h��*���#�1�<�
�>�}�JϮ�H¹��9��h��N���u�u�u�0�$�}�W���Y���F��h_�����4�
�9�
�9�.���Y����l��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	����V9��^ �����&�<�;�%�8�8����T�����1��@���
�<�
�&�>�3����Y�Ƽ�\��DF��Dۊ�
�y�%�d���(����Ƽ�W��h[�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`���&����R��[
��U���;�_�u�u�w�}�W���&�ד�lS��Y1����u�
�d�0�b�W�W���Y�Ʃ�@�N��U���u�u�%�d���(���
���F��_��*ߊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&�ד�lP��G1�����
�<�u�&�>�3�������KǻN��*���0�c�4�
�;���������Z��G��U���'�6�&�}��l��������WJ��h_�����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������1��C���
�9�|�u�?�3�}���Y���F�G1�*���
�%�#�1�>�����DӖ��9��1��*���n�u�u�u�w�8����Y���F�N��*���0�c�4�
�;��������C9��h��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lW��R1�����<�u�&�<�9�-����
���9F���D���c�<�
�<��.����	����	F��X��¥�d�
�
�y�'�l�(���&����F��_��*܊�%�#�1�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	����V9��V�����u�=�;�_�w�}�W���Y�Ƽ�W��hX�����2�i�u�
�f�8�A�ԜY���F��D��U���u�u�u�u�'�l�(���&����Z�
N��Dۊ�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���&����F�	��*���b�a�%�n�]�}�W��	�Փ�lV��G1��ʴ�&�2�u�'�4�.�Y��s���C9��R1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K����^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h\�\���=�;�_�u�w�}�W���Y����V9��V�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s�����h��U��2�%�3�
�f��E�ԜY�Ƽ� 9��^��Hʧ�2�b�d�_�w�}�Z���&����V��G1��ʴ�&�2�u�'�4�.�Y��s���C9��R1�*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ԓ�@��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӖ��l��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&����V��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�G1����u�h�3�
���8���K¹��T9��X����u�x�%�f�2�l�(�������@��YN�����&�u�x�u�w�-�D���H¹��l��h�����%�:�u�u�%�>����	������D�����
��&�g��.�(��s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�o����K�����YNךU���u�u�u�u���(�������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�f�2�l�(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�J����F���*��n�_�u�u�z�-�D���H����l�������%�:�0�&�w�p�W���	�Փ�lW��V�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�E݁�
����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���K����lT��G�����_�u�u�u�w�}�W���&����l��A��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�-�D���H����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����lU��h_�I����;�1�
�2�0�#�������V6��h��*���
�`�g�_�w�}�Z���&����U��G1��ʴ�&�2�u�'�4�.�Y��s���C9��R1�*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ԓ�@��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӖ��l��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&����U��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�G1����u�h�6�
���6�������lU��R1�����d�d�n�_�w�}�ZϮ�J����9��h��U���<�;�%�:�2�.�W��Y����lU��h_�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K����^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h\�\���=�;�_�u�w�}�W���Y����V9��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�J����9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ي�
�
�%�#�3�<����Y����V��C�U���%�f�0�d�6�����
����l��TN����0�&�4�
�2�}��������B9��h��G���8�g�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�}����s���F�N�����0�d�4�
�;�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�G1�����4�
�9�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�
�
�
�w�`��������9��dךU���x�%�f�0�e�<�(���Y����T��E�����x�_�u�u���(݁�	����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�g�
�&��l�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�g�1�0�E���PӒ��]FǻN��U���u�u�
�
���������R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�n���E�ƪ�l��u�����'�2�d�g�l�W�W���TӖ��l��h�����4�&�2�u�%�>���T���F��1��F���
�9�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��_��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���u�=�;�_�w�}�W���Y�Ƽ� 9��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&���� 9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��h]��*���h�3�
�����������U��=d��U���u�
�
�
��-��������]F��X�����x�u�u�%�d�8�C���&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�g�3�8�e�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��F���Y����l�N��U���u�%�f�0�c�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�f�0�a�4��1�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u���(���DӅ��]	��h�����&�4�0��9�/����Hù��T9��V����u�x�%�f�2�h�����ƭ�@�������{�x�_�u�w��(���&����_��D�����:�u�u�'�4�.�_�������C9��P1������&�g�
�$��F�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�e�;���P����[��=N��U���u�u�u�
���(������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�
�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�-�D���O���P
��X
�����
�4�6�1�3�2����&����l��h_�F�ߠu�u�x�u���(ف�	������^	�����0�&�u�x�w�}�����Г�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!�e�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���F��R ��U���u�u�u�u�'�n��������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�f�2�k���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W���&����[��[1�����0�8��&�6�8�4�������l^��R	��C��_�u�u�x�w��(���&����_��D��ʥ�:�0�&�u�z�}�WϮ�J����l��A�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�o����K��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�E݁�
����O�C��U���u�u�u�u�w�-�D���N����E
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�%�d�8�@���&����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���&����F������
�0�8��$�<��������l��h��*��f�_�u�u�z�}�(܁�&˹��l�������%�:�0�&�w�p�W���	�Փ�l^��G1�����&�2�
�'�4�g��������C9��N��*���
�&�$���)�E�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����W�N�����u�u�u�u�w�}�����ޓ�C9��SN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�'�n��������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����V9��S�����c�n�_�u�w�p�����ߓ�C9��SN�����u�'�6�&�y�p�}���Y����V9��V�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�E݁�
����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���K����lT��G�����_�u�u�u�w�}�W���&����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w��(���&����_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
��-��������T9��D��*���6�o�%�:�2�.�����֓�C9��SB��*ފ�
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�����4�
�9�|�w�5��ԜY���F�N��A���e�4�
�9��3����E�Ƽ�9��1��*���n�u�u�u�w�8����Y���F�N��*ފ�
�
�%�#�3�4�(���Y����lR��h^�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l��h�����4�&�2�u�%�>���T���F��1��E���
�<�
�&�>�3����Y�Ƽ�\��DF��A���e�u�
�
������Y����V9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(ہ�&ù��l��R�����0�e�_�u�w�}�W������F�N��Uʥ�a�0�e�<��4�W��	�ғ�lV��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(ށ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��1��*���
�;�&�2�6�.���������T��]���
�
�
�%�!�9�W���&����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�C���H����E
��N�����u�u�u�u�w�}�����ד�C9��S1��*���u�h�%�a�2�l������ƹF�N�����_�u�u�u�w�}�W���&����R��[
�����2�i�u�
���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
������Ӈ��Z��G�����u�x�u�u�'�i��������T9��D��*���6�o�%�:�2�.�������C9��R1�����y�%�a�0�f�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��A���d�4�
�9�~�}����s���F�N�����0�d�<�
�>�}�JϮ�M����l�N��Uʰ�&�u�u�u�w�}�W���	�ғ�lW��Y1����u�
�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�a�2�o��������l��h�����%�:�u�u�%�>����&ǹ��9��h��Yʥ�a�0�g�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ފ�
�
�%�#�3�t����Y���F�N��U���
�
�
�%�!�9���������h��*���#�1�_�u�w�}�W������F�N��Uʥ�a�0�g�4��1�(���
���F��1��G���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��R1�����<�u�&�<�9�-����
���9F���*���
�;�&�2�6�.���������T��]���
�
�y�%�c�8�E�������lR��h\�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`�����ԓ�C9��SG�����u�u�u�u�w�}�WϮ�M����l��D��I���
�
�
�n�w�}�W�������9F�N��U���u�
�
�
��3����E�Ƽ�9��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�C���J����E
��^ �����&�<�;�%�8�8����T�����h��*���#�1�<�
�>���������PF��G�����%�a�0�f�6����	�ғ�lU��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&ǹ�� 9��h��*���&�2�i�u���(܁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ғ�lU��G1�����
�<�u�h�'�i��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�c�8�D���&����R��P �����&�{�x�_�w�}�(ہ�&����l��h�����%�:�u�u�%�>����&ǹ�� J��hZ��*ي�'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����V9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���u�h�%�a�2�n����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ފ�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(ہ�	����l��D�����2�
�'�6�m�-����
ۖ��l��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�a�0�a�4��1�^������F�N��U���%�a�0�a�6���������Z�G1�����4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hZ��*ފ�;�&�2�4�$�:�W�������K��N�����0�a�<�
�>���������PF��G�����%�a�0�a�w��(���&����F��1��A���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ǹ��9��h��\���=�;�_�u�w�}�W���Y����V9��^ �����h�%�a�0�c�W�W���Y�Ʃ�@�N��U���u�u�%�a�2�i���������h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R��[
�����2�4�&�2�w�/����W���F�G1�����4�
�9�
�9�.����
����C��T�����&�}�
�
�������Ƽ�9��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ғ�lS��G1�����!�0�u�u�w�}�W���YӖ��l��h�����<�
�<�u�j�-�C���L����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���
�;�&�2�k�}�(ہ�&ƹ��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�M����l��D�����2�
�'�6�m�-����
ۖ��l��N��A���`�%�0�y�'�i��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�a�0�`�6�����Y����l�N��U���u�%�a�0�b�4�(���Y����lR��h[�U���u�u�0�&�w�}�W���Y�����h��*���&�2�i�u���(ځ�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�a�0�c�4��1�(���
����@��YN�����&�u�x�u�w�-�C���O����E
��^ �����&�<�;�%�8�}�W�������C9��R1�����9�y�%�a�2�k��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
��-����PӒ��]FǻN��U���u�u�
�
����������@��S��*ފ�
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�a�2�k��������l��R�����0�c�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��A���c�<�
�<�w�.����	����@�CךU���
�
�
�
�9�.����
����C��T�����&�}�
�
��q�����Г�A����*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l��h�����|�!�0�u�w�}�W���Y����lR��hX�����2�i�u�
���L���Y�����RNךU���u�u�u�u���(ف�����Z�G1�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ғ�lQ��G1�����
�<�u�&�>�3�������KǻN��*ފ�
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�c�8�@���&������h��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9�� 1��*���|�u�=�;�]�}�W���Y���C9��R1�����9�
�;�&�0�a�W���&����R��[
�U���u�u�0�&�w�}�W���Y�����h��*���#�1�<�
�>�}�JϮ�M����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p�����ѓ�]9��PN�����u�'�6�&�y�p�}���Y����V9��^ �����&�<�;�%�8�}�W�������C9��R1�U���
�
�
�'�0�}�(ہ�&Ĺ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
����������[��=N��U���u�u�u�
���(���
���F��1��B�ߊu�u�u�u�;�8�}���Y���F�G1�����<�
�<�u�j�-�C���N����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��h[��*ڊ�%�#�1�u���(߁�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�`�2�m�������G��d��U���u�u�u�%�b�8�G���&����Z��^	��Hʥ�`�0�e�4��1�L���Y�����RNךU���u�u�u�u���(߁�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�`�0�g�4�(���&����T��E��Oʥ�:�0�&�%�b�8�G���&ƹ��9��R	����0�e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��R1�����9�|�u�=�9�W�W���Y���F��1��E���
�<�u�h�'�h���s���F�R��U���u�u�u�u�w�-�B���I����@��S��*ߊ�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�`�0�d�4��1�(���
����@��Y1�����u�'�6�&���(���&����_�G1�����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h��*���#�1�|�!�2�}�W���Y���F��h[��*ۊ�%�#�1�<��4�W��	�ӓ�lW��G1���ߊu�u�u�u�;�8�}���Y���F�G1�����4�
�9�
�9�.���Y����V9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ƹ��9��h��U���<�;�%�:�2�.�W��Y����lS��h_�����2�4�&�2��/���	����@��h[��*���%�`�0�d�'�8�[Ϯ�L����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�b�8�F���&����F��R ��U���u�u�u�u�'�h��������TF���*���n�u�u�u�w�8����Y���F�N��*ߊ�
�
�;�&�0�a�W���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�`�2�o��������l�������%�:�0�&�w�p�W���	�ӓ�lT��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��@���g�4�
�9�{�-�B���K����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(݁�	����O��_�����u�u�u�u�w��(���&����_��Y1����u�
�
�
��-����s���F�R��U���u�u�u�u�w�-�B���K����E
��^ �����h�%�`�0�e�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�`�0�g�>�����
������T��[���_�u�u�
���(���
����@��Y1�����u�'�6�&���(���UӖ��l��h�����
�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h[��*؊�%�#�1�|�#�8�W���Y���F���*���
�;�&�2�k�}�(ځ�&��ƹF�N�����_�u�u�u�w�}�W���&����Z��^	��Hʥ�`�0�g�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
��-��������T9��D��*���6�o�%�:�2�.�����Փ�C9��SB��*ߊ�
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�����4�
�9�|�w�5��ԜY���F�N��@���f�4�
�9��3����E�Ƽ�9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�
�
�%�#�3�4�(���Y����lS��h]�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l��h�����4�&�2�u�%�>���T���F��1��F���
�<�
�&�>�3����Y�Ƽ�\��DF��@���f�u�
�
������Y����V9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(ځ�&����l��R�����0�f�_�u�w�}�W������F�N��Uʥ�`�0�f�<��4�W��	�ӓ�lU��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(ہ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��1��*���
�;�&�2�6�.���������T��]���
�
�
�%�!�9�W���&����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�B���M����E
��N�����u�u�u�u�w�}�����ғ�C9��S1��*���u�h�%�`�2�i������ƹF�N�����_�u�u�u�w�}�W���&����R��[
�����2�i�u�
���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
������Ӈ��Z��G�����u�x�u�u�'�h��������T9��D��*���6�o�%�:�2�.�������C9��R1�����y�%�`�0�c�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��@���a�4�
�9�~�}����s���F�N�����0�a�<�
�>�}�JϮ�L����l�N��Uʰ�&�u�u�u�w�}�W���	�ӓ�lR��Y1����u�
�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�`�2�h��������l��h�����%�:�u�u�%�>����&ƹ��9��h��Yʥ�`�0�`�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ߊ�
�
�%�#�3�t����Y���F�N��U���
�
�
�%�!�9���������h��*���#�1�_�u�w�}�W������F�N��Uʥ�`�0�`�4��1�(���
���F��1��@���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��R1�����<�u�&�<�9�-����
���9F���*���
�;�&�2�6�.���������T��]���
�
�y�%�b�8�B�������lS��h[�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`�����ӓ�C9��SG�����u�u�u�u�w�}�WϮ�L����l��D��I���
�
�
�n�w�}�W�������9F�N��U���u�
�
�
��3����E�Ƽ�9��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�B���O����E
��^ �����&�<�;�%�8�8����T�����h��*���#�1�<�
�>���������PF��G�����%�`�0�c�6����	�ӓ�lP��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&ƹ��9��h��*���&�2�i�u���(ف�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ӓ�lP��G1�����
�<�u�h�'�h��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�b�8�A���&����R��P �����&�{�x�_�w�}�(ځ�&Ź��l��h�����%�:�u�u�%�>����&ƹ��J��h[��*܊�'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����V9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���u�h�%�`�2�k����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ߊ�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(؁�	����l��D�����2�
�'�6�m�-����
ۖ��l��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�`�0�b�4��1�^������F�N��U���%�`�0�b�6���������Z�G1�����4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h[��*݊�;�&�2�4�$�:�W�������K��N�����0�b�<�
�>���������PF��G�����%�`�0�b�w��(���&����F��1��B���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ƹ��9��h��\���=�;�_�u�w�}�W���Y����V9��^ �����h�%�`�0�`�W�W���Y�Ʃ�@�N��U���u�u�%�`�2�j���������h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R��[
�����2�4�&�2�w�/����W���F�G1�����4�
�9�
�9�.����
����C��T�����&�}�
�
�������Ƽ�9��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ӓ�l^��G1�����!�0�u�u�w�}�W���YӖ��l��h�����<�
�<�u�j�-�B���A����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���
�;�&�2�k�}�(ځ�&˹��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L����l��D�����2�
�'�6�m�-����
ۖ��l��N��@���m�%�0�y�'�h��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�`�0�m�6�����Y����l�N��U���u�%�`�0�o�4�(���Y����lS��hV�U���u�u�0�&�w�}�W���Y�����h��*���&�2�i�u���(ׁ�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�`�0�l�4��1�(���
����@��YN�����&�u�x�u�w�-�B���@����E
��^ �����&�<�;�%�8�}�W�������C9��R1�����9�y�%�`�2�d��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
��-����PӒ��]FǻN��U���u�u�
�
����������@��S��*ߊ�
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�`�2�d��������l��R�����0�l�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��@���l�<�
�<�w�.����	����@�CךU���
�
�
�
�9�.����
����C��T�����&�}�
�
��q�����ߓ�A����*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l��h�����|�!�0�u�w�}�W���Y����lS��hW�����2�i�u�
���L���Y�����RNךU���u�u�u�u���(ց�����Z�G1�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�Г�lV��G1�����
�<�u�&�>�3�������KǻN��*܊�
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�a�8�G���&������h��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��1��*���|�u�=�;�]�}�W���Y���C9��R1�����9�
�;�&�0�a�W���&����R��[
�U���u�u�0�&�w�}�W���Y�����h��*���#�1�<�
�>�}�JϮ�O����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p�����֓�]9��PN�����u�'�6�&�y�p�}���Y����V9��^ �����&�<�;�%�8�}�W�������C9��R1�U���
�
�
�'�0�}�(ف�&ù��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
����������[��=N��U���u�u�u�
���(���
���F��1��E�ߊu�u�u�u�;�8�}���Y���F�G1�����<�
�<�u�j�-�A���I����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��hX��*ۊ�%�#�1�u���(ށ�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�c�2�l�������G��d��U���u�u�u�%�a�8�F���&����Z��^	��Hʥ�c�0�d�4��1�L���Y�����RNךU���u�u�u�u���(ށ�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�c�0�f�4�(���&����T��E��Oʥ�:�0�&�%�a�8�F���&Ź��9��R	����0�d�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��R1�����9�|�u�=�9�W�W���Y���F��1��D���
�<�u�h�'�k���s���F�R��U���u�u�u�u�w�-�A���H����@��S��*܊�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�b�0�e�4��1�(���
����@��Y1�����u�'�6�&���(���&����_�G1�����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h��*���#�1�|�!�2�}�W���Y���F��hY��*ڊ�%�#�1�<��4�W��	�ѓ�lV��G1���ߊu�u�u�u�;�8�}���Y���F�G1�����4�
�9�
�9�.���Y����V9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&Ĺ��9��h��U���<�;�%�:�2�.�W��Y����lQ��h^�����2�4�&�2��/���	����@��hY��*���%�b�0�e�'�8�[Ϯ�N����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`�8�G���&����F��R ��U���u�u�u�u�'�j��������TF���*���n�u�u�u�w�8����Y���F�N��*݊�
�
�;�&�0�a�W���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�b�2�l��������l�������%�:�0�&�w�p�W���	�ѓ�lW��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��B���d�4�
�9�{�-�@���H����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(ށ�	����O��_�����u�u�u�u�w��(���&����_��Y1����u�
�
�
��-����s���F�R��U���u�u�u�u�w�-�@���H����E
��^ �����h�%�b�0�f�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�b�0�d�>�����
������T��[���_�u�u�
���(���
����@��Y1�����u�'�6�&���(���UӖ��l��h�����
�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��*ۊ�%�#�1�|�#�8�W���Y���F���*���
�;�&�2�k�}�(؁�&��ƹF�N�����_�u�u�u�w�}�W���&����Z��^	��Hʥ�b�0�d�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
��-��������T9��D��*���6�o�%�:�2�.�����ԓ�C9��SB��*݊�
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�����4�
�9�|�w�5��ԜY���F�N��B���g�4�
�9��3����E�Ƽ�9��1��*���n�u�u�u�w�8����Y���F�N��*݊�
�
�%�#�3�4�(���Y����lQ��h\�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l��h�����4�&�2�u�%�>���T���F�� 1��G���
�<�
�&�>�3����Y�Ƽ�\��DF��B���g�u�
�
������Y����V9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(؁�&����l��R�����0�g�_�u�w�}�W������F�N��Uʥ�b�0�g�<��4�W��	�ѓ�lT��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(܁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��1��*���
�;�&�2�6�.���������T��]���
�
�
�%�!�9�W���&����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�@���J����E
��N�����u�u�u�u�w�}�����Փ�C9��S1��*���u�h�%�b�2�n������ƹF�N�����_�u�u�u�w�}�W���&����R��[
�����2�i�u�
���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
������Ӈ��Z��G�����u�x�u�u�'�j��������T9��D��*���6�o�%�:�2�.�������C9��R1�����y�%�b�0�d�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��B���f�4�
�9�~�}����s���F�N�����0�f�<�
�>�}�JϮ�N����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�lU��Y1����u�
�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�b�2�i��������l��h�����%�:�u�u�%�>����&Ĺ��9��h��Yʥ�b�0�a�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�
�
�%�#�3�t����Y���F�N��U���
�
�
�%�!�9���������h��*���#�1�_�u�w�}�W������F�N��Uʥ�b�0�a�4��1�(���
���F�� 1��A���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��R1�����<�u�&�<�9�-����
���9F���*���
�;�&�2�6�.���������T��]���
�
�y�%�`�8�C�������lQ��hZ�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`�����ғ�C9��SG�����u�u�u�u�w�}�WϮ�N����l��D��I���
�
�
�n�w�}�W�������9F�N��U���u�
�
�
��3����E�Ƽ�9��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�@���L����E
��^ �����&�<�;�%�8�8����T�����h��*���#�1�<�
�>���������PF��G�����%�b�0�`�6����	�ѓ�lS��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&Ĺ��9��h��*���&�2�i�u���(ځ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�lS��G1�����
�<�u�h�'�j��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�`�8�B���&����R��P �����&�{�x�_�w�}�(؁�&ƹ��l��h�����%�:�u�u�%�>����&Ĺ��J��hY��*ߊ�'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����V9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���u�h�%�b�2�h����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(ف�	����l��D�����2�
�'�6�m�-����
ۖ��l��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�b�0�c�4��1�^������F�N��U���%�b�0�c�6���������Z�G1�����4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��*܊�;�&�2�4�$�:�W�������K��N�����0�c�<�
�>���������PF��G�����%�b�0�c�w��(���&����F�� 1��C���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��9��h��\���=�;�_�u�w�}�W���Y����V9��^ �����h�%�b�0�a�W�W���Y�Ʃ�@�N��U���u�u�%�b�2�k���������h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R��[
�����2�4�&�2�w�/����W���F�G1�����4�
�9�
�9�.����
����C��T�����&�}�
�
�������Ƽ�9�� 1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ѓ�lQ��G1�����!�0�u�u�w�}�W���YӖ��l��h�����<�
�<�u�j�-�@���N����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9�� 1��*���
�;�&�2�k�}�(؁�&Ĺ��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�N����l��D�����2�
�'�6�m�-����
ۖ��l��N��B���b�%�0�y�'�j��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b�0�b�6�����Y����l�N��U���u�%�b�0�`�4�(���Y����lQ��hY�U���u�u�0�&�w�}�W���Y�����h��*���&�2�i�u���(؁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�b�0�m�4��1�(���
����@��YN�����&�u�x�u�w�-�@���A����E
��^ �����&�<�;�%�8�}�W�������C9��R1�����9�y�%�b�2�e��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
��-����PӒ��]FǻN��U���u�u�
�
����������@��S��*݊�
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�b�2�e��������l��R�����0�m�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���m�<�
�<�w�.����	����@�CךU���
�
�
�
�9�.����
����C��T�����&�}�
�
��q�����ޓ�A����*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l��h�����|�!�0�u�w�}�W���Y����lQ��hV�����2�i�u�
���L���Y�����RNךU���u�u�u�u���(ׁ�����Z�G1�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�l_��G1�����
�<�u�&�>�3�������KǻN��*݊�
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�`�8�N���&������h��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��1��*���|�u�=�;�]�}�W���Y���C9��R1�����9�
�;�&�0�a�W���&����R��[
�U���u�u�0�&�w�}�W���Y�����h��*���#�1�<�
�>�}�JϮ�N����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p�����ߓ�]9��PN�����u�'�6�&�y�p�}���Y����V9��^ �����&�<�;�%�8�}�W�������C9��R1�U���
�
�
�'�0�}�(؁�&ʹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
����������[��=N��U���u�u�u�
���(���
���F�� 1��L�ߊu�u�u�u�;�8�}���Y���F�G1�����<�
�<�u�j�-�@���@����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��hW��*ڊ�%�#�1�u���(߁�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�l�2�m�������G��d��U���u�u�u�%�n�8�G���&����Z��^	��Hʥ�l�0�e�4��1�L���Y�����RNךU���u�u�u�u���(߁�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�l�0�g�4�(���&����T��E��Oʥ�:�0�&�%�n�8�G���&ʹ��9��R	����0�e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��R1�����9�|�u�=�9�W�W���Y���F��1��E���
�<�u�h�'�d���s���F�R��U���u�u�u�u�w�-�N���I����@��S��*ӊ�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�
9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�l�0�d�4��1�(���
����@��Y1�����u�'�6�&���(���&����_�G1�����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h��*���#�1�|�!�2�}�W���Y���F��hW��*ۊ�%�#�1�<��4�W��	�ߓ�lW��G1���ߊu�u�u�u�;�8�}���Y���F�G1�����4�
�9�
�9�.���Y����V9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ʹ��9��h��U���<�;�%�:�2�.�W��Y����l_��h_�����2�4�&�2��/���	����@��hW��*���%�l�0�d�'�8�[Ϯ�@����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�n�8�F���&����F��R ��U���u�u�u�u�'�d��������TF���*���n�u�u�u�w�8����Y���F�N��*ӊ�
�
�;�&�0�a�W���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%��&�9��i����N����Z������,� �
�b�1��Eځ�H����W	��C��D���u�8�
�c�>�;�(��&���9F������!�a�
� �f�d�(��E����C9��Y����
�u�u�:���G���&����l��d��Uʥ��&�9�
�a�;�(��K����[�Q=��4����!�d�
��(�F��&���F��@ ��U��u�u�8�
�a�4�(���H����CU�=N��U���0� �!�&�1��Gځ�J�����T�����d�
�u�u�8��(���A�ߓ�O��N�����g�<�<�<�g�>��������F9��V��F��u�u�u�u�w�<�(���
����S��^�����}�8�
�
���@���&����l��G��U��|�0�&�u�w�}�W�������]��[�*��n�u�u�'�#�o��������G9��D�� ��l�%�u�h�]�}�W���Y����\��h��@���e�"�0�u�#�-�D�������F9��1��]���h�r�r�u�;�8�}���Y���R��X ��*���`�d�e�_�w�}����&����l ��^�*��i�u�u�u�w�}��������_��hZ�Eʢ�0�u�!�%�d�4����&����U��G\��\��r�r�u�9�2�W�W���Y�ƭ�l��D�����a�e�n�u�w�/��������F9��1��U��_�u�u�u�w�-��������9��^�����}�8�
�
���(���A�ߓ�N��S��D���0�&�u�u�w�}�WϿ�&����G9��[��A��_�u�u�0��0�F���&����Q��G\��H���8�
�
�
�a�;�(��K����K	��V�����
�#�
�|�]�}�W���&����l��B1�@���u�h�}�8���(�������l��O�����:�&�
�#��t�}���Y����G��h�����e�e�%�u�j�u����&����Z_��B1�@؊�g�4�1�&�;�)�ށ�J����V��h�N���u�&�9�!�'��(���A�ד�F�F�����<�<�<�3��k�(������V
��Z�����
�m�
�g�l�}�Wϭ�����9��h��D��
�g�i�u�f�}����Q����~3�� ����
�;�3��'��(���H����CU������!�9�d�
�c�m�W�������l�N�����%�
�
� �n�d����D������YN��&��� ��;� ��n����	����l ��W�����u�%�6�;�#�1�Fځ�M���V
��L�N���u�&�9�!�'��F���&����l��S��D���=�;�}��/��#ݰ�����l��Q�����
� �d�m��n�JϿ�&����G9��[��E���0�&�u�e�l�}�Wϭ�����9��Q��Lߊ�g�i�u�d�w�5����*����2��x��Gي�;�3��%��(�O���	���R��X ��*���`�a�e�u�;�8�U���s���@��C��*���3�
�d�e�'�}�J�������CP��1��*��m�%�u�'�$�1����&�ד�F9��Z��G��u�u�&�9�#�-�(�������9��R��]���
�8�c�<�1��Oց�KӉ��@��C��*��� �l�`�%�~�W�W�������C9��h��D��
�f�i�u�w�}�W�������l��1��*��a�%�u�=�9�u����&����l ��^�*��e�u�u�d�~�8����Y���F��G1�����9�d�
�e�l�}�Wϭ�����l��B1�B���u�h�_�u�w�}�W���&����Z9��hV�*��"�0�u�!�'�4�������� 9��^��H��r�u�9�0�]�}�W���Y����\��h��@��e�_�u�u�:��(���&�ѓ�F9��V��G��u�d�u�=�9�u����&�ד�F9��V��D��4�
�:�&��+�D��Y����D��d��Uʡ�%�f�<�<�>�;�(��&���F�N�����9�6��d��(�O���	���R��X ��*���f�e�u�9�2��U�ԜY�Ƹ�C9��h�����d�a�%�u�j��Uϩ�����Z��SF��*����g��!�e�����	����l ��_�*��u�u�<�;�3�<�(���
����^��G�����w�w�_�u�w�0�(�������
T��G\��H���w�"�0�u�$�:����*����2��x��Gي�;�0�%��f�;�(��&���F��P ��]���6�;�!�9�f��^������D��N�����`�
�d�3��l�C���Y���G��_�� ��a�
�f�s�'�m�G߁�&�ד�F9��X��F��u�u�!�%�b��(���@�ӓ� F�F����
� �l�b�'�}�W���K�֓�l��B1�B���|�_�u�u�:��(���@�ӓ� F�d��U���u�4�
�:�$��ׁ�?ӑ��]F��Z��*���l�l�%�}�~�`�P���Y����l�N��Uʴ�
�:�&�
�!��L���YӒ��lS��h��L���
�e�g�%�w�`�U�������
��h8��E���
�e�m�%�w�}��������E^��qG�����w�w�_�u�w�0�(ځ�&����U��]��G��u�d�u�=�9�u����&����_��N�����:�&�
�#���W�������l�N�����3�
�d�a�'�}�J�ԜY���F��h�����#�
��"�2�}����¹��lW��1��]���h�r�r�u�;�8�}���Y���R��X ��*���
�n�u�u�#�-�@ց�����l��S��U���u�u�!�%�b�;�(��&����[����*��� �l�d�%��t�J���^�Ʃ�@�N��U���!�%�l�
�"�d�D���B�����hV�����d�e�%�u�j�u����H����W��h����8�
�`�<��(�F��&���9F���*���3�
�d�c�'�}�J�ԜY���F��G1�����d�a�%�u�?�3�_���&�֓�F9��^��G��u�u�d�|�2�.�W���Y�����hW�����d�g�%�n�w�}����@ƹ��l_��h�I����-� ��9�(�(�������C9��1��*��
�g�m�x�f�9� ���Y����F�C��L݊� �d�a�
�f�a�W���������C1�*���0�%��f�1��F���	����F��S�����|�_�u�u�:��F���&����l��S��D���=�;�}�<�9�9����4����])��h\�����-�
�
�
�"�l�G݁�K���@��R
�����;�!�9�d���^ϻ�
���]ǻN�����
� �l�l�'�}�J���[ӑ��]F��^	��³�
���g��)�E܁�����l0��h��L���%�|�k�&�0�8�_�������l
��1��\���9�0�w�w�]�}�W���&����ZP��B1�F؊�g�i�u�d�w�5��������V��B1�DҊ�a�h�4�
�8�.�(���&����_��^�����u�8�
�
�����J����[�L�����}�:�
�
�"�e�N���Y�ƭ�l��D��Ҋ�|�0�&�u�g�f�W�������l ��]�����h�}�8�
��(�N���	�ƣ���h[�����
�g�
�g�l�8�ϼ�����