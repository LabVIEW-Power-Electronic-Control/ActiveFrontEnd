-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�8����_��1��F���
�
�l�f�%�0����Y����V��^��U���u�u�u�u�:�0����Y�����^ ��O���7�:�>�n�]�}�W���Y���W��C��U���u�;�0�0�w�`�D��s���F�N�����!�u�u�u�w�3����Y���FǻN��U���u�u�0�
�>�8�W���Y����T��S�����u�n�_�u�w�2����Y���F������u�u�u�;�$�9��������G	��V�����u�:�;�:�g�f�}���Y���F��N��U���o�<�u�!��2���s���F�N��U���u�u�o�:�#�.��������V��EF�����x�u�:�;�8�m�L���Y���F��S
��U���u�u�;�&�3�1��������AN��^
��X���:�;�:�e�l�W�W���Y���P��N��U��<�u�!�
�8�4�L�ԜY���F�S_��U���u�o�<�u�#�����&����\��@����1�"�!�u�~�}�W���Y�����N��U���u�;�&�1�;�:����Y���F���U���u�u�o�<�w�)�(�����ƹF�N�����;�<�,�u�]�<��������VF��[N��U���c�`�d�3�g�;�D���&����U��V���ߠ&�2�4�u�3�/�(���Y�ƿ�W9��P�����:�}�"�1�?�l��������F��N�����4�'�,�<�w�/����IӒ��^��D��X���:�u�!�
�8�4�(������W��C��U���;�:�e�n�]�5��������Q
��E��Oʸ�8�4�'�,�m�}�������\��E��R��|�_�4�!�>�(�ϭ�����@��RN����;�n�_�!�%�?���� ����^��[��ʧ�8�o�#�'�6�1�W���[����X9��ZL����<� �0�'�:�.����Cӕ��Z��=�����!�u�4�
�#�1�W��������^��ʼ�u�0�
�,�2�W��������v7��a/��;���������!���Cӕ��Z��=d�����_�_�0�:�.�<����&����W9�������u�4�1�e�w�?����Y�����E^�����h�4�1�e�]�p��������G��D�����3�u�u�u�>�}�4���&����t#��V
��E���u�0�
�<�2�l�W������F�N�����e�!�%�i�w�2����Y���A�=N��U���9�0�_�u�w�}�W�������l��R�����e�_�u�u�w�3�W���s�˿�]��D�����&�4�0�:�]�3�W�������9l��Z�����6�0�&�e�w�/����Yۅ��F�U���ߊu�u�3�}�;�z����Y����P
��
N��R���=�;�u�u�w�}�������A��N�����u�u�u�u�w�}����DӔ��%��a1��!����4�1�e�#�-�^���Y���F��Y
���ߊu�u�;�u�1�W��������@]Ǒ=�����,�4�6�&��g�������P
��N�����u�u�u�<�w�>�Ȼ�����]��[��U��|�!�0�_�w�}�W����ί�F�_��U���;�_�u�u�w�}�W����λ�F�_��U���;�_�u�u�w�}�W���Y�ƾ�^N��y8��;����}�1�'�~�}�JϺ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���_�;�u�'�4�.�L�Զ����G
��=d�����,���n�"�8�>���W����_	��T1�C���9�n�_�;�>�$�ߟ�N����U9��Q1�����
�l�f�<�]�}�W�������l�N��Uʑ�!��1�=�m��#���+��� T��N��U����1�0�&�6�:�W���7����aF��\�U���u�u��1�2�.����Y�ƅ�g#��eN�U���_�u�u�:�#�u�W���Y����V��T��;ʆ�����]�}�W���Y����	F��=��*����n�u�u�w�}��������	F��=��*����
��������
����[F�N��"���u�|�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�&�}�W���Y����)��t1��6���}�4�4�<�#�}�W���6����V�=N��U���u�1�'�&�f�g�>���-����t/��a+��:���1�'�&��3�5�Z��=����|F��d��U���u�6�d�o��}�#���6����9F�N��U���u�u�����0���s���F�S_��U���������4���Q����d��_N�Dʑ���u�|�l�8�ϻ�����9l��T�����'�u�'�=�8�}�G��L����lV��h]�����d�`�u�&�w�}����������Y�Dӳ�e�3�f�3���N�������@l�N��Uʥ�'�u�_�u�w�}�W���Y����	F��=��*����n�u�u�w�}�W�������\��yN��1��������f�W���Y���F��R^��U��������W�W���Y���F��T�� ����
�����#���s���F�N�����d�o��u���8���&����|4��N��U���u�u�6�d�m��W���&����p]ǻN��U���u�u�d�o��}�#���6����e#��x<�U���u�u�u�u� �l�Mϗ�Y����)��tG�U���0�1�6�8�8�8��Զs����ZǻN��E��`�d�3�e�1�n����&����l��h;��Uʶ�8�:�0�!�:��@��@����U9��Q��*��f�'�8�u�w�-�������F�N�����h�u�9�y�w�}�W�������[�V
�����y�u�u�u�w�>�G��Y����9F�N��U��h�u�e�_�w�}�W�������X��S
����_�u�u�u�w�8�W�������F�N�����k�1�y�u�w�}�Wϩ�H���D��d�����'�=�!�6�"�8�}��