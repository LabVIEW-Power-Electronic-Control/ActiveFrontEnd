-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�8����_��1��F���3�f�g�f���(���Y���F�P�����_�u�u�u�w�}�W���&����F�N�����u�h�w�9�4��W���Y���F�
�����u�u�o�<�#�:���Y���F�N��U���4�<�!�u�w�}�W�������	[�NךU���u�u�u�u�2�����Y����Z��P��O���_�u�u�n�]�}�W�����ƹF�N��U���'�u�u�u�w�3��������l��C�����!�x�u�:�9�2�G��s���F�N��E���u�u�o�<�w�)�(������F�N��Uʤ�u�u�u�u�m�2�ϭ�����Z��R��±�<�!�x�u�8�3���B���F�N�����u�u�u�u�9�.��������V��EF�����x�u�:�;�8�m�L�ԜY���F�T�U���u�o�<�u�#�����B���F�N�����u�u�u�o�>�}��������E��X�����=�d�1�"�#�}�^���Y���F���U���u�u�u�;�$�9������ƹF�N��U��u�u�u�u�w�(�W���&����P9��T��]���1�=�d�1� �)�W���s���F�N�����u�u�u�u�9�.�������F�U�����0�!�!�n�]�W��������A��C��ʸ��b�d�l���(܁�����_��h��*���u�&�_�&�0�<�W���ù��CF��D�����6�#�6�:��*����Hӂ��]��G����;�9�4�1�f�)���
����\��h�����4�<�!�x�w�2����I���G����*���4�u�&�4�%�$�_���Ӌ��l��RC�U���&�1�9�2�4�+����Yۂ��W��N�����u�|�u�&�6�8�W���������T�����'�4�n�_�#�/����Y����A��C��U���!�<�2�u�6�)����ӕ��l��D��ʺ�u�4�u�u�6�4��������_	��h��W���!�'�7�!�w�<�(�������@��Y	����<� �0�'�:�.�����ƾ�^F��A�����u�&�8�8�#�-�L������G��f;��4���������2���8����@��Y	����<�u�_�8�:�/�(�������F��h^����0�&�}�1�%�t�}������F�V
��E���%�i�u�1�%�f�Z­�����Z��E�����
�3�_�u�w�}����6����}2��r<�����|�k�8�8�$�'�Z�������F�N��U���1�'�
�8�w�`�_������F�G�U���u�0�&�u�w�}�W���Y�ƭ�W��C��I���1�'�n�u�w�}������ƴ��C�����'�;�9�!��3����	����@��=�����,�4�6�&��g�������P
��N�����u�u�u�<�w�>�Ȼ�����]��[��U��|�!�0�_�w�}�W����ί�F�_��U���;�_�u�u�w�}�W���I���A��t!��*�����}�1�%�����B���F�N��ʼ�n�u�u�0�3�4�L��Ӗ��P��d�����,�4�6�&��(����CӖ��P��F����u�7�2�;�w�}�WϿ��ד�^�
N����_�x�,�!�2�4�W�������V9��Qd��U���<�u�����2���Q����O���*���0�d�u�=�9�}�W���Y���R��1����u�:�=�'�w�c�P���B���F��[�����u�u�u�u�6�9�F���	���R��UךU���u�;�u�3�]�p��������G��D�����_�;�u�'�4�.�L���&����A��T����u�'�6�&�w�>����s����]FǻN�����9�r�#�;�w�3�W���Y���O��_��U���u�u�<�u�4�l�J���^�Ƹ�V�N��U���u�u�<�u� �l�J���^�Ƹ�V�N��U���u�u�u�u�%�0�4���&����t#��V
��D���%�|�o�u�f�}�W���Y���F��Y
���ߊu�u�u�u�w�}�F��Y����p)��h'��0���}�1�'�
�:�t�L�ԜY���F��SN��N���u�0�1�<�l�8�Ϯ�����lǑR �����_�_�<�'�%�}�2���s����z#����*���<�
�d�a�6�1�}������^V�� [�L���
�
�
� ���N�������@l�N�����6�}�u�u�w�}�3���.����\��y:��0���h�d�_�u�w�}�W�������R��T��;����u�h�a�]�}�W���Y����V��^
��U������u�j�o�L���YӖ��GF�N��U���'�&�!�o��}�#���6����9F�N��U���u�u�����0���s���F�V
�����u�u�����0���/����aN��S�����!�u�u�u���8��B���F���U���������}���Y���BV�!��U���
���
��	�%ǚ�����G�_��:����e�n�u�w�}�WϿ�����F��~ ��!�����
����6�������W��N�1����u�|�_�w�}�W�������z(��c*��:���n�u�u�u�w�*�F��0�Ɵ�w9��p'�����u�u�u�d�m��W���&����p9��t:��]���4�<�!�u�w�}�8���6���9F�N��U��o������0���/����aN��C�����x�d����}�^������]��NUװ���<�0�!�'�w�/�ϱ�Y�֍�S����*���
� �
�
�n�l������F��Z�����8��b�d�n��(���&���� 9��_��*ڊ�4�u�&�u�w�}�WϮ����F�N��U���6�>�o��w�	�(���0��ƹF�N��U���1�'�u�u���3���>����v%��eUךU���u�u�u�u�2�}�W���*����|!��d��U���u�u�u�$�w�}�"���-����t/��a+��:��u�u�u�u�w�}����H����}F��s1��2������n�w�}�W���Y����VW�'��&������_�w�}�W���Y�ƨ�\��yN��1��������f�W���Y���F��R_��U��������W�W���Y���F��T�� ����
�����#���B����������;�n�_�_�2�4�}���Y�֍�S����*���
� �
�
�n�l��������\�T�����!�8��b�f�d�(߁�&����U9��W�*���
�4�_�u�w�2�ϳ�	��ƹF�N�����k�6�>�_�w�}�W�������X��S
����_�u�u�u�w�8�W�������F�N�����k�$�y�u�w�}�WϿ����F��S�����u�u�u�u�4�l�J�����ƹF�N��D��u�d�_�u�w�}�W���Y����VW�N��U���$�u�k�$�~�W��������G��B����