-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��b�d�l���(�����A�=N��U���6�>�o��w�	�(���0��ƹF��G1�����u��
���L���YӇ��@��CN�<����
���l�}�WϿ�&����\��b:��!�����n�u�w�<�(�������f2��c*��:���n�u�u�4��8����Y����`2��{!��6�ߊu�u�;�-�g�g�>���-����t/��a+��:���f�u�:�;�8�m�L���YӇ��A��E ��U��� �u��
���(���-��� W��X����n�u�u�4��8����H����f2��c*��:���
�����l��������l�N��*���o��u����>���B����lǑV�����!�'�u�0�6�}�ϳ�8����_��1��D���&�_�u�u�8�.��������]��[����o������M���H��ƹF��X �����4�
�:�&��2����Y�Ɵ�w9��p'��O���e�n�u�u�4�3����Y����g9��1����o������!���6�����Y��E���h�w�e�e�f�f�W�������R��V��!���g�3�8�d�m��3���>����v%��eN��U���;�:�e�u�j��G��I��ƹF��X �����4�
��&�d�;���Cӵ��l*��~-��0����}�u�:�9�2�G���D����W��UךU���:�&�4�!�6��#���M����lU�=��*����
����u�W������F��L�D��w�_�u�u�8�.��������l��h��*���u��
����2���+����W	��C��\��u�e�e�e�u�W�W�������]��G1��*���
�&�
�u�w�	�(���0����p2��F����!�u�|�o�w�l�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�F��Cӵ��l*��~-��0����}�u�:�9�2�G���D����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>�������� F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EW��T��!�����
����_�������V�S��E��u�u�6�;�#�3�W�������l
��1��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�e�n�u�w�>�����ƭ�l��D�����f�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��d�d�d�w�]�}�W���
������T�����`�
�u�u���8���&����|4�]�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��1�Oʆ�������8���O�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��1�F��������4���Y����W	��C��\��u�e�e�e�f�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�e�G��*����|!��h8��!���}�u�:�;�8�m�W��[����V��UךU���:�&�4�!�6�����&����l ��T��!�����
����_������\F��T��W��d�d�d�e�f�f�W�������R��V�����
�#�g��m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����W��d��Uʶ�;�!�;�u�'�>�������� P�=��*����
����u�FϺ�����O�
N��E��e�d�d�e�l�}�WϽ�����GF��h�����#�c���w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��H����W��_�W�ߊu�u�:�&�6�)��������_��h^��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�1��Cӵ��l*��~-��0����}�d�1� �)�W���C���W��_�E��n�u�u�6�9�)����	����@��A_��D���u��
����2���+������Y��E���h�w�e�e�g�l�G��B�����D��ʴ�
�:�&�
�!�o�1���Cӵ��l*��~-��0����}�d�1� �)�W���C���W��_�D��n�u�u�6�9�)����	����@��A_��F���u��
����2���+������Y��E���h�w�e�e�g�l�F��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���`�1�"�!�w�t�M���I����D��N�����!�;�u�%�4�3����O����	F��s1��2������u�b�9� ���Y���F�^�E��u�u�6�;�#�3�W�������l
��1��3�������w�}�#���6����e#��x<��@���:�;�:�e�w�`�U��H����W��_�D��d�d�d�d�f�l�F��H����W��_�D��d�n�u�u�4�3����Y����\��h��G��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�e�n�u�w�>�����ƭ�l��D������o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�d�d�n�w�}��������R��X ��*���d�d�o����0���/����aF�N�����u�|�o�u�g�m�G��I���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>�����ӓ�\��c*��:���
�����}�������	[�^�E��u�u�6�;�#�3�W�������l
��1�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����b��u�u���8���&����|4�[�����:�e�u�h�u�l�F��H����W��UךU���:�&�4�!�6�����&����l^��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�o�D��*����|!��h8��!���}�u�:�;�8�m�W��[���9F������!�4�
�:�$�����I����g"��x)��*�����}�f�3�*����P���V��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��I���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����W��UךU���:�&�4�!�6�����&����F��d:��9�������w�n��������\�^�E��u�u�6�;�#�3�W�������l
��1�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*۔�o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�d�w�]�}�W���
������T�����g�e�o����0���/����aF�
�����e�u�h�w�g�f�W�������R��V�����
�#�g�d�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�m�U�ԜY�Ư�]��Y�����;�!�9�`�f�}�W���&����p9��t:��U��1�"�!�u�~�g�W��I���9F������!�4�
�:�$��݁�Y�Ɵ�w9��p'��#����u�d�1� �)�W���C���D��N�����!�;�u�%�4�3����L����	F��s1��2������u�c�9� ���Y���F�_�W�ߊu�u�:�&�6�)��������_��h_�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��A]��D���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��d�w�_�u�w�2����Ӈ��P	��C1��Gߊ�u�u��
���(���-���R��X����u�h�w�e�g�m�G��I����V��^�D��u�u�6�;�#�3�W�������l
��hY�Oʆ�������8���Nӂ��]��G��H���d�d�e�d�l�}�WϽ�����GF��h�����#�d�e�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�f�
��m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�d�f�m�L�ԜY�ƿ�T����6���&�u�u����>���<����N��S�����|�o�u�e�g�m�U�ԜY�ƭ�G��B�����0�6�1�;�w�}�������F��C�� ���3�8�0�6�3�3�W�������l ��T�����9�<�u�;�9��}���Y����R
��G1�����0�
��&�f�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�6����&����V��T��!�����
����_������\F��d��Uʦ�2�4�u�4�%�l���Cӵ��l*��~-�U���&�2�4�u�6�/�F���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����
�
�1�'�$�l�Mύ�=����z%��r-��'���e�1�"�!�w�t�}���Y����R
��V��D���d�o�����4�ԜY�ƿ�T�������$�u�u����>���<����N��
�����e�n�u�u�$�:��������l��E��E��������4���Y����W	��C��\�ߊu�u�<�;�;�6����&����	F��s1��2���_�u�u�<�9�1����&����\��c*��:���
�����h��������l�N�����u�4�'�g�6�9����Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����
�
�0�u�w�	�(���0��ƹF��^	��ʾ�'�
�
�d�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������^��1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������9��P1�G���u��
����2���+������Y��E��u�u�&�2�6�}�(���K�ԓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����K����lT��N�&���������W��Y����G	�UךU���<�;�9�$��(�C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���'�2�g�f�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������l ��\�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�/����K����	F��s1��2������u�g�9� ���Y����F�D�����8�
�c�3��n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
�0�
�g�g�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���`�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�_9��G]�����g�`�o����0���/����aF�N�����u�|�_�u�w�4����
����^��Q��Bۊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l��h\�E��������4���Y����\��XN�N���u�&�2�4�w�8�(���M����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)�ہ�����S�=��*����
����u�W������]ǻN�����9�!�%�f��(�A���	����`2��{!��6�����u�`�3�*����P���F��P ��U���
�b�'�2�e�k�W���-����t/��a+��:���`�1�"�!�w�t�}���Y����R
��G1�����0�
��&�e�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�.��������lT��N�&���������W������\F��d��Uʦ�2�4�u�%�$�:����&����GU��D��U����
���l�}�Wϭ�����R��^	�����e�u�u����L���Yӕ��]��G1��؊�f�'�2�g�n�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���
�g�m�o���;���:����g)��^�����:�e�n�u�w�.����Y����@��Y1�����b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����@��Y1�����g�e�u�u���8���&����|4�N�����u�|�_�u�w�4����
����Z��h��*��l�o�����4���:����V��X����n�u�u�&�0�<�W����ԓ�9��P1�D���u��
����2���+������Y��E��u�u�&�2�6�}����H����lT��N�&���������W������\F��d��Uʦ�2�4�u�7�6�.����&���� V��N�&���������W������\F��d��Uʦ�2�4�u�7�6�.����&����U��T��!�����
����_�������V�=N��U���;�9�!�%�>�;�(��K����	F��s1��2������u�g�9� ���Y����F�D�����8�
�
�0��n�D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1����Lǹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Bہ����� ^�=��*����
����u�W������]ǻN�����9�;�8�0��?�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u� �5�/����/����lT��N�&���������W��Y����G	�UךU���<�;�9�!�'�4�E܁�����9��T��!�����
����_�������V�=N��U���;�9�!�%�>�o�(���&����\��c*��:���
�����}�������9F������;�8�0�
�2�9��������U��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�3����&����a	��S��#���2�g�`�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��l��Q��G���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����A��]�U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Aׁ�����9��T��!�����
����_�������V�=N��U���;�9�!�%�a�����J���5��h"��<������}�w�2����I��ƹF��^	��ʻ�8�0�
�7���(���H����CU�=��*����
����u�BϺ�����O��N�����4�u� �7�%�<����L����lT��N�&���������W��Y����G	�UךU���<�;�9�!�'�4�(�������R��N�&���������W������\F��d��Uʦ�2�4�u�8��l�Eہ�����V�=��*����
����u�W������]ǻN�����9�;�8�0��8��������e9��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����]��e������d�'�2�e�e�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h^�D���<�3�
�a�a�-�W���-����t/��a+��:���a�1�"�!�w�t�}���Y����R
��h^�D���<�'�2�g�n�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������D�����
��&�`�1�0�C��*����|!��d��Uʦ�2�4�u�%�$�:����H���$��{+��N���u�&�2�4�w��B���K����F9��Z��G��������4���Y����\��XN�N���u�&�2�4�w��B���K����V��W�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��8����K����A��Z�U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������V��N��1��������}�E�������V�=N��U���;�9�%�e�o��(������� P��N�&���������W������\F��d��Uʦ�2�4�u�
�b�l�D���&����R��T��!�����
����_�������V�=N��U���;�9�%�e�`��(�������R��N�&���������W������\F��d��Uʦ�2�4�u�
�b�j�E���&����R��T��!�����
����_�������V�=N��U���;�9�%��$�1�(�������lT�� N�&���������W��Y����G	�UךU���<�;�9�!�'�o�(���&����\��c*��:���
�����o��������l�N�����u�8�
�
��(�A���	����`2��{!��6�����u�c�w�2����I��ƹF��^	��ʡ�%�c�<�3��h�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V��*���<�;�3�
�d��G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������f�
� �g�`�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��؊�d�3�
�f��l�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��1�����l�
�d�o���;���:����g)��\����!�u�|�_�w�}����Ӗ��R
��V�� ��d�%�u�u���8���&����|4�X�����:�e�n�u�w�.����Y����_T��1��*��
�d�o����0���/����aF�
�����e�n�u�u�$�:����&����T��B1�F���u�u��
���(���-���U��X����n�u�u�&�0�<�W�������F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�%�(���&����lT��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�#�-�O���&����CW�=��*����
����u�FϺ�����O��N�����4�u�8�
�"�o�N���Y�Ɵ�w9��p'��#����u�`�u�8�3���B�����Y�����&�9�
�f�1��O؁�H����g"��x)��*�����}�f�3�*����P���F��P ��U���0�
� �g�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��V ��*ۊ� �g�d�%�w�}�#���6����e#��x<��@���:�;�:�e�l�}�Wϭ�����G��1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������l ��Y�����u��
����2���+������Y��E��u�u�&�2�6�}�E���&����CT�=��*����
����u�FϺ�����O��N�����4�u�8�
�f�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʼ�8�
� �f�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��*���f�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��Q��Fӊ�g�o�����4���:����W��S�����|�_�u�u�>�3�ϭ�&����U��[��F��������4���Y����W	��C��\�ߊu�u�<�;�;�0��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��m����N����\��c*��:���
�����}�������9F������&�
�8�
�6�)����L����\��c*��:���
�����l��������l�N�����u�8�
�
�"�n�N���Y�Ɵ�w9��p'��#����u�`�u�8�3���B�����Y�����c�3�
�l��o�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��Z��A���
�c�
�d�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������^��1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������9��hZ�*��o������!���6���F��@ ��U���_�u�u�<�9�1����N���� P��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���J�ߓ�F��d:��9�������w�l�W������]ǻN�����9�%�&�3��m�(��Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V�����`�3�
�f��o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��D���&�
� �a�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��Dي� �a�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������l ��Y�����u��
����2���+������Y��E��u�u�&�2�6�}����I����^��G_��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�l�(���M�ѓ�F��d:��9�������w�m��������l�N�����u�
�%�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �a�f�'�}�W���&����p9��t:��U���1�"�!�u�~�W�W���������h]�����e�
�d�o���;���:����g)��[����!�u�|�_�w�}����Ӓ��lU��Q��Eߊ�g�o�����4���:����S��S�����|�_�u�u�>�3�Ϫ�	����U��_��G��������4���Y����W	��C��\�ߊu�u�<�;�;�-�%�������U��Y��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����S��N�&���������W������\F��d��Uʦ�2�4�u�8��d����K����\��c*��:���
�����}�������9F������!�%�d�3��m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����3�
�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���`�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CP��R�����3�
�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���`�`�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��]�����2�;�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��^��A���
�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����U��[��G��������4���Y����\��XN�N���u�&�2�4�w�?��������U��W��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�D���&����CT�=��*����
����u�BϺ�����O��N�����4�u�0�
�:�e����H����\��c*��:���
�����h��������l�N�����u�-�
�0�:���������Z��1�����d�
�f�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lP��^1��*��
�a�o����0���/����aF�
�����e�n�u�u�$�:����5����V9��E��Dڊ�
�4�!�3��n�(��Cӵ��l*��~-��0����}�e�1� �)�W���s���@��V��9������!�%��N���&����CT�=��*����
����u�GϺ�����O��N�����4�u�8�
�g�4����O¹��\��c*��:���
�����k��������l�N�����u�8�
�d�>�;�(��&���5��h"��<������}�a�9� ���Y����F�D�����8�
�g�<�1��@ځ�H����g"��x)��*�����}�c�3�*����P���F��P ��U���
�f�<�3��j�(��Cӵ��l*��~-��0����}�c�1� �)�W���s���@��V��*��� �c�l�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��[\��D���
�f�
�g�m��3���>����v%��eN��Gʱ�"�!�u�|�]�}�W�������^��1��*��
�d�o����0���/����aF�
�����e�n�u�u�$�:��������l �� \�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�/�F���&����CT�=��*����
����u�W������]ǻN�����9�'�<�<�>�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʤ�<�
� �b�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��U1�����
�
� �b�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h8��G��
� �c�l�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*��� �b�b�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����A9��1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4����	����9��h��G���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l �� V�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����
V��N�&���������W������\F��d��Uʦ�2�4�u�
��(�@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�d�<�3��d�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
� �b�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V�����
� �m�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V��Aڊ� �b�g�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����G��^��*���m�e�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��h]�����`�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lT��^1��*��
�d�o����0���/����aF� N�����u�|�_�u�w�4��������9��Q��Gڊ�d�o�����4���:����W��S�����|�_�u�u�>�3�Ϭ�/�Փ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�$�<�����K����	F��s1��2������u�g�9� ���Y����F�D�����
�4�g�a��(�O���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʡ�%�f�
�
�"�e�E���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����f�
�
� �o�e����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��#��
� �m�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���l�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��G9��Q��Dڊ�d�o�����4���:����V��X����n�u�u�&�0�<�W���&�ޓ�l ��]�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K����U��W��G��������4���Y����W	��C��\�ߊu�u�<�;�;�3� �������U��Z��F��������4���Y����\��XN�N���u�&�2�4�w�0�(�������
S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�6�%�$����L˹��\��c*��:���
�����}�������9F������!�%�f�
��(�N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0� �!�;�#�4����Nƹ��\��c*��:���
�����}�������9F������!�%�f�
��(�N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���:�
�
�
�"�d�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�
�
�
�"�d�A���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����0�
�;�&�1��Aׁ�J����g"��x)��*�����}�u�8�3���B�����Y�����'�0�e�1�:�/����&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�9�:��������9��T��!�����
����_�������V�=N��U���;�9�7�8�%�8�G�������V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�9�8����&����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�:�2�;��������9��T��!�����
����_�������V�=N��U���;�9�;�2�$�>��������V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:�l����I�ޓ�F��d:��9�������w�m��������l�N�����u�'�0�2���(�������9��T��!�����
����_�������V�=N��U���;�9�7�8�%�8����&����l��N��1��������}�GϺ�����O��N�����4�u�
�4�e�l�(���&����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w���������V��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�#�-�C݁�&����Q��G_��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u��<�E��&����Q��G\��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u�2�.�����ד�F9��\��F��������4���Y����\��XN�N���u�&�2�4�w�0�(�������V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�/�(ށ�����9��T��!�����
����_�������V�=N��U���;�9�!�%�c��(���H����CT�=��*����
����u�W������]ǻN�����9�%��&�;��(���&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�B߁�&����W��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%�9�)�ށ�&����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�7�:�/����&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�3�1��������9��h_�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��X�����
�
� �d�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Y�����d�3�
�d�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E����
�d�<�3��l�E���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�:�
�
�"�l�Bׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����3�:�
�
�"�l�C߁�K����g"��x)��*�����}�u�8�3���B�����Y�����&�6�f�;�#�4����H�֓�F��d:��9�������w�m��������l�N�����u�8�g�3��l�A���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�
�
�d�>�;�(��M����	F��s1��2������u�g�9� ���Y����F�D�����'�0�2�d�>�;�(��K����	F��s1��2������u�g�9� ���Y����F�D�����
�4�g�d��(�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�F�������
P��N�&���������W��Y����G	�UךU���<�;�9�3�'�3��������_��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������A9��D1��D���
�g�c�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��D��*���3�
�g�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[�����g�c�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӏ��l��R1�����d�
�
� �f�m�(��Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V�� ���'�4�&��d�;�(��I����	F��s1��2������u�f�}�������9F������%��&�9��o����K�ғ�F��d:��9�������w�j��������l�N�����u�8�
�f�1��D���	����`2��{!��6�����u�d�3�*����P���F��P ��U���
�
� �d�e��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������!�g�
� �f�o�(��Cӵ��l*��~-��0����}�l�1� �)�W���s���@��V��*���d�3�
�f�c�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��؊�d�3�
�f�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����
�a�<�3��n�E���Y�Ɵ�w9��p'��#����u�f�1� �)�W���s���@��V��*���
� �d�c��i�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��h8��G��
�
�4�!�4�.�(���H����CU�=��*����
����u�W������]ǻN�����9�!�%�`�����O����\��c*��:���
�����}�������9F������%��&�9��h����J�ԓ�F��d:��9�������w�i��������l�N�����u�
�
�g�1��D���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ��9�
�
�"�l�G߁�J����g"��x)��*�����}�l�3�*����P���F��P ��U���0� �!�d�����I˹��\��c*��:���
�����}�������9F������'��c�3��i�C���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�g�3��n�E���Y�Ɵ�w9��p'��#����u�a�1� �)�W���s���@��V�����g�<�3�
�c�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������!�g�
� �f�n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��#��
� �d�f��l�Mύ�=����z%��r-��'���l�1�"�!�w�t�}���Y����R
��h8��G���3�
�a�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��a1�����a�g�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��h[�����a�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lS��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�+����G9��h��D��
�a�o����0���/����aF�
�����e�n�u�u�$�:����&����l ��Z�*��o������!���6���
F��@ ��U���_�u�u�<�9�1��������l ��[�*��o������!���6���
F��@ ��U���_�u�u�<�9�1��������\%��C�����&��3�
�b�i����Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T����*���3�
�`�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������hX�����`�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��D���
�g�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�C���u�u��
���(���-���S��X����n�u�u�&�0�<�W�������lT��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l��B1�D؊�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�ғ�l ��[�*��o������!���6�����Y��E��u�u�&�2�6�}�����ד�l ��[�*��o������!���6�����Y��E��u�u�&�2�6�}����L����F9��V��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:�n����L�Г�F��d:��9�������w�m��������l�N�����u�0�
�8�e�4����L�ғ�F��d:��9�������w�m��������l�N�����u�0�
�8�b�4����O�ԓ�F��d:��9�������w�m��������l�N�����u�8�
�m�>�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�
��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�
��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʻ�!�&�9�!�'��(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�n����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�(�������9��T��!�����
����_�������V�=N��U���;�9�'��o�;�(��N����	F��s1��2������u�d�}�������9F������%��&�9��o����O�֓� F��d:��9�������w�n�W������]ǻN�����9�'��d��(�F��&���5��h"��<������}�n�9� ���Y����F�D�����
�4�g�c��(�F��&���5��h"��<������}�n�9� ���Y����F�D�����
�0� �!�e��(���H����CR�=��*����
����u�W������]ǻN�����9�'��l�1��@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ��9�
�a�>�>��������F9�� V��F��������4���Y����\��XN�N���u�&�2�4�w�0�(�������Q��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��8����J����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�%��Fف�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�A���&����l��N��1��������}�D�������V�=N��U���;�9�%��$�1�(�������Q��h�Oʆ�������8���Hӂ��]��G�U���&�2�4�u���(���H����CR�=��*����
����u�@Ϻ�����O��N�����4�u�
�4�e�k�(���H����CU�=��*����
����u�W������]ǻN�����9�!�%�c�����L˹��\��c*��:���
�����}�������9F������%��&�9��i����N�ޓ�F��d:��9�������w�i��������l�N�����u�
�
�b�1��@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ��9�
�
�"�l�Nف�J����g"��x)��*�����}�l�3�*����P���F��P ��U���
�
� �d�f��C��*����|!��h8��!���}�m�1�"�#�}�^�ԜY�ƿ�T�������c�
� �d�o��D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Bۊ� �d�e�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C9��D��*���3�
�m�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_�����m�g�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��hX�����m�a�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƣ�^��h��6���<�4��!���(���H����CW�=��*����
����u�W������]ǻN�����9�!�%�b��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�b�
� �f�e�(��Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V�����b�3�
�m�g�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��C��BҊ� �d�l�
�e�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������R����
� �d�e��o�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��Z��A���3�
�m�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������hX�����
�m�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z��ۊ� �d�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��X��D���
�m�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^�� 1�����m�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1��*���d�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�CT��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CS��1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������
9��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����l��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��h��D��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������_9��GW��D���
�l�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���3�
�l�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Dڊ�d�3�
�l�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��G1�����0�
��&�a�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������F��u!��0���_�u�u�<�9�1��������F��R�����3�
�e�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��Z��*���;��&�9���(���K����CT�=��*����
����u�CϺ�����O��N�����4�u� �7�%�/��������\��h��G��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������l��B1�D݊�d�o�����4���:����R��X����n�u�u�&�0�<�W�������V��Y	�����0�
�
�
�"�o�Eށ�K����g"��x)��*�����}�u�8�3���B�����Y����m�
�
�
�"�o�Eف�J����g"��x)��*�����}�u�8�3���B�����Y�����c�
�
� �e�n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �g�`��l�Mύ�=����z%��r-��'���g�1�"�!�w�t�}���Y����R
��Z��A���
�e�m�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����C9��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�+����G9��h��G��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	����F
��^�� ��c�
�a�o���;���:����g)��]����!�u�|�_�w�}����ӈ��Q��D	�����
�
� �g�`��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������%�0�<�<�9�;��������l��B1�Aۊ�g�o�����4���:����Q��X����n�u�u�&�0�<�W�������lU��Q��E���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l��B1�Lي�d�o�����4���:����U��S�����|�_�u�u�>�3�ϰ�����A	��S<�� ����g�3�
�f�i����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����
�:�;��$�1�(���&����V��G\��U���
���
��	�%���Mӂ��]��G�U���&�2�4�u�"�?��������V��X��*ۊ� �g�d�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G�� ^��*���g�g�
�d�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƣ�^��h������0�;�0���(���K����CT�=��*����
����u�W������]ǻN�����9�%�e�m���F���&����l��N��1��������}�CϺ�����O��N�����4�u�8�
�f�4����H�ד�F��d:��9�������w�j��������l�N�����u�8�
�d�1��F���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʡ�%�g�
� �e�k�(��Cӵ��l*��~-��0����}�g�1� �)�W���s���@��V��*���3�
�d�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������R����
� �g�`��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h<�� ���f�
� �g�a��C��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�� �����&�9�=�9���(���K����CU�=��*����
����u�FϺ�����O��N�����4�u�<�2�2�-��������_	��h��*���
�
� �g�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1�����
�l�3�
�f�h����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
�
� �g�n��F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������e�l�3�
�g�j����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*���8�
�d�3��o�F���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������3�8�o���;���:����g)��[�����:�e�n�_�w�}��������^V�� [�L���
�%�-�
�e�.�Aہ�Y��ƹF��R �����_�u�u�u�w��Mϗ�-����l�N��Uʛ�����m��#���+���F�N��ڊ���u�u���2��Y���F��X��"����o�����^�ԜY�Ƽ�A�=N��U���u�<�e�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӂ��GF��x;��&���������W��Y����G	�N����u�;�u�:�'�3���s�����G�����e�c�`�d�1�m���&����lW��dd��Uʲ�;�'�6�}�w�}�W���=����Z��T��;����n�u�u�w�}�6�������]��N��!����_�u�u�w�}����
����G�'��0���u�n�u�u�'�/�W�ԜY���F��\N�<����
���l�}�W���YӔ��V�'��&������_�w�}�W�������@V�'��&���������W��Y����G	�UךU���u�u�0�u�w��$���5����l�N��Uʤ�u�u� �u���8���&����|4�[�����:�e�n�u�w�}�WϿ�����F��~ ��!�����
����_������\F��d��U���u�6�d�o��}�#���6����9F�N��U��o������0���/����aF�N�����u�|�|�_�w�}��������V��=dךU���:�%�;�;�w�m�A��Hʀ��l ��1�����u��u�u�0�3����Q���F�*�����!�u�u����L���Y���'��E��'���0�o�����}���Y���r��R�����u�u����}�L���YӖ��GF�N��U���6�>�o��w�	�(���0��ƹF�N�����u�u�����0���s���F�V
�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�&�}�W���Y����)��t1��6���u�d�u�:�9�2�G��Y���F��S
����o��u����>���<����N��
�����e�n�u�u�w�}���Cӯ��`2��{!��6�ߊu�u�u�u�f�g�8���*����|!��h8��!���}�`�1�"�#�}�^���s���V��T�����!�_�_�7�0�3�W�������9��N�����0�!�8��`�l�N���&����l��E1�U���2�;�'�6�:�-�_���Y���"��V9�����k�d�y�u�w�}�Wϟ�����a��RN��U��`�_�u�u�w�}����
����G�	N�\���u�%�'�u�6�}�}���Y���P
��
P�����>�_�u�u�w�}����Y����C9��CBךU���u�u�1�'�$�m�J�������l��E��E�ߊu�u�u�u�2�}�Iϵ�����P��=N��U���u�e�h�u�6�/�F���U���F������d�h�u�4�%�l��������9F�N��U���u�k�>�'�����Y���F��N��U���'�d�$�|�]�}�Wϵ�����fF��T�����!�8��b�f�d�(߁�&�֓�R��d��Uʲ�;�'�6�8�'�u�W���Y����R��^
��U��d�y�u�u�w�}�6�������]��
P��E���_�u�u�u�w�9����.����[�_��U���%�'�u�4�w�W�W���Y�Ư�XF������_�u�u�u�w�8����GӇ��A��=N��U���u�1�'�&�g�`�W����ԓ�W��D����u�u�u�0�w�c����&����JǻN��U���e�h�u�4�%�o���Y���F��S
����h�u�4�'�e�<����
��ƹF�N�����k�>�'�
��8�[���Y�����
P�����g�$�|�_�w�}��������lU��D1�*ۊ�e�o�6�8�8�8�ϳ�8����_��1�����f�;�
�a�f�}�WϹ�������FךU���u�u��h�w�q�W���Y����f+��c/��U��d�_�u�u�w�}����.����[�\�U���u�u�1� ���#���G����9F���ʸ�%�}�u�u�w�}����Y����l��^	�����f�
�e�_�w�}�W������F��V����� �g�f�%�~�W�}�ԶY���F��RN�����!�&�4�0��-�4���
����UF��RN�����8�6�<�0�w�p�W�������l ��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�%��
�$�}�JϿ�&����GW��D��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�_�u�u�w�}�W���Y���F��h-�����i�u�%���.�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h]��\ʡ�0�_�u�u�w�}�W���Y�Ƣ�^��h��*���
�0�
�f�d�a�W�������Q��h[�� ��m�
�f�_�w�}�W���Y���F��Z��*���
�
�0�
�d�i�K�������l��h8�� ��f�
�f�_�w�}�W���Y���F��Z��*���1�:�;�0���(���&����Z�Y�����0�1�:�;�2��(ށ�����9��d��U���u�u�u�u�w�3����&����a	��S��#���2�g�`�u�j�3����&����a	��S��#���
�g�e�%�l�}�W���Y���F���*���'�2�g�f�w�`��������G��h_�*��� �d�c�
�d�l�W������O��N��U���u�u�u�u�#�-�Aׁ�����Q�
N�����1�
�0�8�f�h�!���&����l��[�����:�d�|�_�w�}�W���Y���F��G1��*���'�2�g�m�w�`����¹��l ��]�*��_�u�u�u�w�}�W���Y����ZW��R	��F��i�u�8�
�f�;�(��O����9F�N��U���u�u�u�8���D�������F���*���f�3�
�g�g�-�L���Y���F�N��U���
�
�0�
�d�n�K�������U��_����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C�����;�%�:�0�$�}�Z���YӖ��P��F��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y�����Yd��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ځ�
������F�����
�0�
�f�e�`��������_��G��U���;�u�u�u�w�}�W���YӖ��Q��1��*���
�a�e�i�w��B���K����U��Y����u�u�u�u�w�}�W���	����9��^_�����a�a�i�u��h�F���¹��lW��1��N���u�u�u�u�w�}�WϮ�+����G9��h�����a�b�i�u��<�E��&����R��G]��Aʱ�"�!�u�|�]�}�W���Y���F�C��Gߊ�0�
�a�g�k�}�(���K����U��Z�����f�1�"�!�w�t�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�6�.��������@H�d��Uʥ�:�0�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��|�!�0�_�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C[�����|�4�1�}�:��(���&����[��G1�����9�d�e�|�w�5����Y���F�N��U���`�b�g�<�%�:�E��Y����lV�� 1�����
�c�a�%�l�}�W���Y���F���@���f�<�'�2�e�d�W��	����9��^1��*��c�%�n�u�w�}�W���Y�����R����
�
�0�
�c�i�K���&����lS��Q��@���%�}�a�1� �)�W���s���F�N��U���!�%�g�
�2��C��E�Ƽ�e��h[�����`�a�%�}�d�9� ���Y����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�6�~�<�ϰ��έ�l��E��U���6�;�!�9�0�>�G���PӒ��]l�N��U���u�u�u�%��1�(݁�����S�
N��#���
�
� �a�b�-�L���Y���F�N��U���'�2�g�f�w�`��������l��=N��U���u�u�u�u�w�����K���F��Q��Gӊ�g�_�u�u�w�}�W���Y�ƿ�_9��G]�����g�`�i�u�2���������9��d��U���u�u�u�u�w�.����	ǹ��T9��[��Hʦ�9�!�%�
�"�h�N���B���F�N��U���u�0�
�8�`�/���L�����h��B���
�b�
�g�]�}�W���Y���F�C��G܊�0�
�g�e�k�}����O����T��G_�U���u�u�u�u�w�}����JŹ��T9��^��Hʡ�%�f�
� �b�h���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��F���8�g�|�u�?�3�W���Y���F�N��*���g�a�
�0��o�D��Y���� 9��hV�*��d�u�:�;�8�l�L���Y���F�N��U���4�g�a�
�2��D��E�ƾ�e9��h��M���%�}�c�1� �)�W���s���F�N��U���$�
�&�<�9�j����K����[��U1�����
�
� �m�e�-�L���Y���F�N��U���4�&�2�
��8�(��A���B��D�����3�
�f�
�e�W�W���Y���F�N�����!�d�'�2�e�m�W������9��hV�*��d�u�:�;�8�l�^�ԜY���F�N��Uʦ�2�7�!�'�0�o�O���DӔ��lU��B1�M���}�b�1�"�#�}�@��Y���F�N��U���8�
�c�'�0�o�N���DӔ��lU��B1�M���}�c�1�"�#�}�A��Y���F�N��U���8�
�d�'�0�o�E���DӔ��lW��Q��M܊�g�d�u�:�9�2�F���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�|�#�8�}���Y���F�N�����f�
�0�
�e�m�K�������l ��]����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C�����0�!�&�4�2�u����&����	��C�����0�8�6�<�2�}�Z���YӇ��}5��D�����;�%�:�u�w�/����Yۇ��@��CB�����
�&�y�4��8�}���Y����]l�N��Uʶ�&�u�%���.�W���Y���F�N�����4�
��&�f�;���D��ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u���������T�����2�6�e�|�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��D�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����]��QUךU���u�u�u�u�?�3����-����l ��h_��K�ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�4������E�ƭ�l5��D�����g�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��h��*���k�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=�����3�8�f�_�w�}�W���Y���F��DךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����3�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�`�3�8�c�W�W���Y���F�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!��.�(��Y���F�N��U���;�u�3�_�w�}�W���Y�ƻ�V��G1��*���
�&�
�u�i�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�c�1�0�B�ԜY���F�N��Uʰ�&�_�u�u�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���u�u�;�u�1�W�W���Y���F��R �����
�!�
�&��}�I�ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l����I���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����!�0�&�h�w�W�W���Y���F�N��*���3�8�i�u���/���s���F�R �����n�u�u�0�3�-����
���F��h��F���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�l�(��P����]��Y�����&�3�
�b��l�^�ԜY�ƃ�9��Q��Lފ�d�i�u�!��2����������^�� ���2�0�}�8��j����K����T��UװU���x�u�%�1�9�}����Ӗ��P��N����u�%�1�;��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�%�6�y�6�����
����g9��1�����_�u�u�0�>�W�W���Y�ƥ�N�Y��]���6�;�!�9�0�>�F������R��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�Г�@��G��U���;�_�u�u�w�}�W���	����VF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�8�8�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���Ӈ��Z��G�����u�x�u�u�6���������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�|�w�}�������F���]»�!�}�%�6�9�)���������D�����4�1�}�%�4�3��������[��G1�����0�
��&�f�;���P�Ƹ�V�N��U���u�u�4�
�3�8�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�'�4�,�6�.��������@H�d��Uʴ�
�0�1�
�$�4��������C��R�����0�u�%�&�0�>����-����l ��h[��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\���=�;�_�u�w�}�W���Y����V��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�/����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�<�(�������Z�Q=�����
�
� �g�n��D�ԜY�ƭ�l��B��D��u��!�'�g�l�(���K����CU��=N��U���4�
�<�
�3��G���
������T��[���_�u�u�%�$�:����H�Փ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��]��H���%�6�;�!�;�l�F������l ��\�����:�g�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��G������]F��X�����x�u�u�4��4�(���&����l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�G��u�4�
�:�$��ށ�Y�ƭ�l%��Q��@ʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���NӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�B��u�4�
�:�$��ށ�Y�ƭ�l%��Q��Fʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���LӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�@��u�4�
�:�$��ށ�Y�ƭ�l%��Q��Aʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Z��H���%��
�&��}�������F��h�����#�
�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��BϿ�
����C��R��U���u�u�4�
�>�����L����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������l^��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��D���8�e�4�&�0�����CӖ��P�������7�1�g�|�w�}�������F���]���&�2�7�1�e�t����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l ��h^��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�o����HӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����m�|�u�u�5�:����Y����������7�1�m�|�#�8�W���Y���F������6�0�
��$�o����H���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���K����lW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�f�1�0�EϿ�
����C��R��U���u�u�4�
�>�����*���� 9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��D��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�e�|�!�2�}�W���Y���F��G1�����0�
��&�d�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�a�3�:�n�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�B�ߊu�u�0�<�]�}�W���Y���R��^	�����g�|�!�0�w�}�W���Y�����D�����
��&�a�1�0�D��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�C������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�`�3�8�c�<����Y����V��C�U���4�
�<�
�$�,�$���ƹ��^9��V�����'�6�o�%�8�8�ǿ�&����Q��[����u�0�<�_�w�}�W����έ�l��h��*���|�!�0�u�w�}�W���Y����C9��P1������&�`�3�:�i�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�h����M���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���c�3�8�`�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&����9��D��*���6�o�%�:�2�.��������W9��\��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��D��|�!�0�u�w�}�W���Y����C9��P1������&�c�3�:�h�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�k����L���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}��������Z9��h_�G���u�h�}�8�e�;�(��O����\��E����
�0�:�2�9�4�(�������9��UךU���'�0�2�a��8��������Z9��h_�C���u�h�}�0�$�:����H����V��h����1�9�!�1�8�8�(ށ�����9��UךU���'�0�2�a��8��������l ��^�*��i�u�;�"�>�3��������l��V �����!�1�:�0��(�N���	����F�U�����e�<�
�
�"�l�B݁�K�����R��Aڊ�0�:�2�;�>��(���H����CT��X�����;�!�9�d�f�f�W�������T��h��*���d�d�
�g�k�}��������l��X�����<�3�
�e�o�-�W���Y����\��h��*���_�u�u�'�2�:�(�������W��h�I���;�"�<�;�>��(���H����CU��EN�����<�
�
� �f�o�(��B�����R��*��� �d�a�
�e�a�WǪ�	¹��lW��1��U���7�8�'�0�g�9��������Z9��h_�M���|�_�u�u�%�8����&�ד�l ��_�*��i�u� �1�%�1� �������^��N��U���'�9�"�d�1��F���	����F�U�����<�<�3�
�n��E��Yۈ��@��U�����a�
�f�:�w�����&����l_��h�N���u�7�8�'�2�4��������P��N�U �1�'�9�"�1��G���	�ƣ�	��E�����
�e�g�%�~�W�W�������9��h_�C���u�h�}�8��l����K����R��C��A܊�
� �d�l��o�L���YӅ��A��B1�M���u�h�}�8��k����K����R��C��F؊�
� �l�g�'�t�}���Y����@��h��G���%�u�h�<���L���Yӂ��V��h�����3�
�d�c�'�}�J�ԜY���F��G1�*��� �d�e�
�e�*��������lW��B1�L܊�g�e�u�u�f�t����Y���F������
�
�0�
�d�d�}���Y����G��X ��*���l�m�%�u�j�W�W���Y�Ƹ�C9��h�� ��f�%�u�=�9�u����&����^��F�U���d�|�0�&�w�}�W���Yӕ��]��h��*��`�_�u�u�/�����&����W��N�U���2��3�
�c��F��Y����G	�G�U���3�
�0�8��l����K�ד� F�d��U���u�4�
�:�$�����Iӑ��]F��Z��D���2�g�c�}�~�`�P���Y����l�N��Uʡ�%�b�
�
�"�o�N؁�H���F��h��ڊ�
� �g�l��n�K���Y���F��G1�����9�f�
�u�?�3�_���&����T9��]��\��r�r�u�9�2�W�W���Y�Ƹ�C9��h�� ��l�
�d�_�w�}��������V��_��#���
�g�a�%�w�`�}���Y���C9��[\��M���-�<�3�
�f�e�������Q��E	��*��� �d�m�
�e�m�W���H����_��=N��U���u�
�4�g�f�4����H�Г� ]ǻN�����:�0�!�'��l�(�������9��R�����u�u�u�
�6�o�Fځ�����U��[�����=�;�}�'�2�:�(�������9��^��H��r�u�9�0�]�}�W���Y����_T��h��D���
�f�_�u�w�%�(�������l ��R
�����`��3�
�f��D��Y���F���*���'�2�g�g�w�5��������CR��R	��G���e�u�u�d�~�8����Y���F��R�����3�
�d�
�d�W�W���5����v>��e����
� �c�l�'�}�Jϭ�����Z��R�� �&�2�0�}��3��������V��h�����
�f�
�d�w�}��������C9��Y����
�|�n�u�w�4�(�������^9��1�����
� �c�`�'�}�Jϭ�����Z��R��§�&�/�}�;�>�3�Ǫ�	����Z9��hX�*��y�d�|�_�w�}����&����U��N�U��u�=�;�}�:��G���&����CR������!�9�m�e�w�1����[���F��Z�� ��b�%�u�h�u�� ���Yە��]��C��Dۊ� �f�b�%�~�c�����έ�l��D��Ҋ�|�u�9�0�u��}���Y����l0��B1�@���u�h�1�4�$�:�(���K�Փ�]ǻN�����
� �g�f�'�}�JϷ�����U��[��D��u�:�;�:�a�t�}���Y����lW��S
����i�u�8�
�����J����W�_�����:�e�n�u�w�6����&����V��R�����c�<�3�
�b��F��Y����W	��C��\�ߠu�u�x�u�6�/�F���IӇ��Z��G�����u�x�u�u�<�/�(ށ�ù��@��h����%�:�0�&�6�����	����l��F1��*���
�&�
�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�~�}����s���F�N�����
�
�0�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���X��h_�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���'�d�6�d�6�.��������@H�d��Uʾ�'�
�
�0��.����	����	F��X��´�
�0�u�%�$�:����&����GT��D��\���u�7�2�;�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��D���u�=�;�_�w�}�W���Y�Ƨ�A��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}����H����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�W�������9��S�����h�!�%�g�>�;�(��&���F�N�����u�|�_�u�w�<��������@��S�����
�
� �c�b�-�_��T����\��XN�N�ߊu�u�x�>�%��(���Y����T��E�����x�_�u�u�6�/�E���I����Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=�����3�8�d�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�)����Y���F�N�����g�6�e�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����R��1��E��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����
�
�0�u�$�4�Ϯ�����F�=N��U���'�g�6�d�6�.���������T��]���6�y�4�
�>�����*����9��Z1����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��D��\���!�0�u�u�w�}�W���YӍ��A9��T�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�6����&����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W�������9��h\�*��i�u�!�
�8�4�(�������]��Y�����:�&�
�#�c�m�W�������V��h<�� ���g�
� �g�`�-�^��Y����R��h��G���%�u�h�_�w�}�W�������9��h\�*��"�0�u�<�9�:����L����V�
N��R���9�0�_�u�w�}�W�������lT��Q��M݊�d�_�u�u�2�����&����T��G\��H���<�;�<�
��8�(��@Ӈ����h[�����
�d�m�%�~�W�W�������P9��Y�����
�d�e�%�w�`�_���&����9��h_�A���u�:�u�%�4�3����H���9F� ��*���
� �l�c�'�}�J�������G9��P1�M���;�u�8�
�a�4����Aù��]ǻN�����'�
�:�
��(�F��&���F��R	����� �l�c�%�w�2�W�������l
��h_����u�0�&�2�5�)�F���&����l��S��*���g�a�
� �f�j�(��H�ƨ�D��_�N���u�;�"�<�9�4�(���@�ғ� F������a�
� �l�n�-�_������\F��UךU���:�
�0�
�:�d�ށ�����9��R��W���"�0�u� �$�:����&����lU��1��*��c�%�|�k�"�.����Q����\��h��*��|�0�&�u�g�f�W�������V
��Z�����
�c�c�%�w�`�U���������^	��¥�e�m�
�
��(�F��&���F��D�����%�6�;�!�;�h�F���Y����D��d��Uʻ�8�0�
�7���(���H����CT�
N�����2�6�#�6�8�u��������C9��Y����
�|�x� �$�:��������W��R��D����3�
�e�a�-�^��Y����F��E1�����f�3�
�g�g�-�W��
����\��h����� �&�2�0��-��������9��C�����;�1�3�%�9�9�(�������l0��B1�Eފ�f�|�_�u�w�(��������lS��B1�M܊�f�i�u�u�w�}�Wϰ�����R��a1�����g�e�%�u�?�3�_���&�ޓ�F9�� \��F��u�u�d�|�2�.�W���Y��� ��h �����'�
�d�
��(�F��&����F�Y�����7�
�
� �f�n�(��E��ƹF�N�� ���'�4�&��f�;�(��O����D��F�����
� �d�d��n�G���Y�����RNךU���u�u�-�
�8�8����&����e9��h_�C���n�u�u�;�:�8�(�������]��S��#���3�
�e�d�'�}�Jϭ�����Z��R�� �&�2�0�}��h�F�������lT��G��U���<�;�1�!�'�h�(�������9��G�U���;�8�0�
�2�9��������K9�� 1��*��`�%�u�h�$�9��������G	��B �����}�
�`�d�d�4�(���&����F�B �����}�8�
�e�>�;�(��H����]ǻN�� ���'�;�0��"�9����H����U��h�I���d�u�=�;��0�(�������V��N�����:�&�
�#��t����Y���9F� �����;�0�� �3�9�!���&����l��S��D���=�;�}�8��d����K�Г�F�V�����
�#�
�|�2�.�W��B�����U�����1�#�'�9� ��F���&����l��S�� ���'�'� �1�2�(����L����W��h�G���:�;�:�g�~�W�W�������l��Y
�����:�
�
� �e�m�(��E�Ƣ�^��h�����&�9�
�
��(�E��&���F��@ ��U��n�u�u�;�:�8�(�������F
��a1�����d�a�%�u�j�.��������V��EF�����}�;�<�;�3�-�%�������l��R	��A��y�`�|�_�w�}��������]��D��*���
� �g�e��o�K�������T��A�����;�<�;�1�9�0��������V��C1�����e�e�%�|�|�(�����έ�l��D�����d�|�_�u�w�(��������a��[��*ߊ� �g�e�
�e�a�W���&����P9��T��]���<�;�1�;�:�8�(�������F
��a1�����d�a�%�|�|�(�����έ�l��D�����d�|�_�u�w�(��������a��[��*���g�e�
�d�k�}��������E��X�����0� �&�2�2�u�(�������9��E��G��|�g�|�n�w�}��������_5��[��*݊� �g�b�
�d�a�W���Y�����R����
� �g�`��n� ���Yۖ��9��h\�C���}�|�h�r�p�}����s���F�G1�����
�m�3�
�f�e���Y����F��E1�����9�
�
� �e�j�(��E��ƹF�N��*��� �!�g�
�"�o�C؁�Jӑ��]F��h�� ��f�
�g�e�w�}�F�������9F�N��U���0� �!�f��(�E��&����F�Y�����"��<�<�6�����&¹��lW��1��U��%��9�
�b�;�(��M����F�N�����u�|�_�u�w�(��������Z��V�����
� �d�g��l�K���&����lS��Q��@���%�}�u�u�w�2����I��ƹF��A�����d�3�
�d�g�-�W��Q����A��^_��*���d�f�
�g�6�9����M˹��U��^�����_�u�u�#�%�1� ���&����l��S�����'�0�<�<�1��Nف�KӇ����h]�����
�c�
�g�l�}�WϮ�I����9��h��D��
�g�i�u�$�1����J����U��X�����'�&�9�!�'�m�ށ�����9��UךU���
�`�b�g�>�;�(��M����[�D�����f�<�3�
�a�e����ӕ��l��^��*���d�g�
�g�l�}�WϮ�I���� 9��h��D��
�f�i�u�w�}�W���	����F
��[�� ��g�
�a�"�2�}����N¹��lW��1��]���h�r�r�u�;�8�}���Y���C9��[\��F���
�b�m�%�l�}�WϮ�I���� 9��Q��A���%�u�h�_�w�}�W���&����_�� 1��*��c�%�u�=�9�u����N����R��h�E���u�d�|�0�$�}�W���Y����l0��1�*���d�a�
�f�]�}�W���L�ד�l��Q��D���%�u�h�_�w�}�W�������l
��S��:���;�0�
�
��(�E��&����[����@���g�<�
�0��i�G��Y���O��[�����u�u�u�
�b�l�D���&����R��d��Uʥ�e�m�
�
��(�E��&���FǻN��U��� �7�'�9�6�4����0����l0��h��G��
�g�"�0�w�-�G��&����A��]�]���h�r�r�u�;�8�}���Y���C9��_��*���0�
�f�d�]�}�W�������lW��^1��*��g�%�u�h�'��݁�H����U��h�F���:�;�:�g�~�W�W���&����_��1�����a�m�%�u�j�-�!���&ǹ��lW��1��]��1�"�!�u�a�f�W���	����F
��]�� ��b�%�u�h�$�9��������G	��E�����;�<�;�1�#�-����Nʹ��J��G�U���%��&�9��i����J�֓� F�F�����
�7�
�
�2��D��_Ӈ��P	��C1��Gފ�|�_�u�u�w�}����
����S��B1�M؊�a�%�:�u�w�/����Q����_T��1�����
�4�!�3��n�O���P�����^ ךU���u�u�
�0�"�)�Eځ�����9��R�����9�
�c�<�4�.�(�������U��h����u�u�u�
�2�(���&���� ^��GZ��\��u�%�6�;�#�1�F��I��ƹF��Y
�����&�n�_�u�w���������Z9��h_�G���u�h�%��;��F���&����l��_�����:�g�|�_�w�}�W���	����F
��X�� ��f�
�a�%�8�}�W�������C9��[\��G���
�f�g�%�~�}�Wϼ���ƹF�N��*��� �!�g�
�"�l�Dׁ�M���C9��[\��G���
�f�g�%�l�}�W���YӖ��V��C1�*���d�f�
�a�f�}�JϿ�&����G9��1�E��u�u�0�1�'�2����s���l�N��'���9�
�b�3��i�A���&����\��E�����
�4�g�`��(�F��&���F�U�����u�u�u�%��.����N����R��h�I���
�4�g�`��(�F��&����F�N�����&�9�
�b�1��C���	����Z�V�����
�#�
�}�~�W�W����Ƽ�\��DUװU���%��&�9��j����&����l��S��*���g�c�3�
�`�m����Nӂ��]��X����u�
�0� �#�o�(���H����CT�
N�� ���'�4�&��%�:�E��Y����G��Z�� ��`�
�g�n�w�}����
����_��B1�A݊�f�i�u�!�'�h�(���&����@��G1�����9�f�
�|�]�}�W�������lU��Q��E���%�u�h�}�#�-�Bہ����� ^������!�9�m�e�w�}����M����V��h�N���u�%��&�;��F���&����l��S�����0�
�2��2�1�!���&����l��_�����:�f�|�s�$�3��������Z	��Q�����%��<�3��m�F���Y�Ƣ�^��h��&���9��3�
�g�n����Kӂ��]��G����u�
�0� �#�n�(���H����CU�
N�� ���'�4�&��b�/���N���R��X ��*���a�e�n�u�w�W�W���&����_��1��*��g�%�
�'�4�g��������l0��1�*���4�!�6�&��(�F��&���F�U�����u�u�u�%��.����J����Q��h�I���
�4�g�g����������U��Y����u�u�u�u�'�����&�Փ�F9��\��A��u�h�4�
�8�.�(���&����l�N��ʥ�:�0�&�_�w�}�}���Y����@��h]�����b�m�%�
�%�>�MϮ�������V��C؊� �d�f�
�d�W�W�������F�N�����&�9�
�a�1��@���	�����V��C؊� �d�f�
�d�W�W���Y�Ƽ�a��[��A���
�b�m�%��t�K���	����@��A_��]���_�u�u�;�w�/����B���FǻN��*��� �!�f�
�"�l�Eف�M����PF��G�����%��9�
�d�;�(��A����9F����ߊu�u�u�u��8����Jƹ��lW��1��U��%��9�
�d�;�(��A����9F�N��U���0� �!�f��(�F��&���F������!�9�d�d�g�f�W�������A	��D����u�
�0� �#�n�(���H����CT�
N�� ���'�4�&��b�/���N�ƭ�WF��G1�*���d�l�
�g�l�}�WϮ�+����G9��h��G���
�f�i�u�#�-�Aׁ�����Q������!�9�f�
�~�W�W���&����_��1��*��m�%�u�h��)���&����U��H�����;�!�9�m�g�}�W���&�ѓ�F9��\��F��u�u�%��$�1�(�������S��N�U»�8�0�
�2��8����N����W��h�F���:�;�:�f�~�{��������V��^�����!�0�%��>�l����H�ӓ�F�Y�����2��0�9��j����H�ѓ� N��
�����e�|�_�u�w������Г�\��h��D��
�g�i�u�#�-�Bށ�����T��X�����;�!�9�d�f�f�W���	����F
��^_�� ��a�
�a�i�w�(��������l ��\�*��d�u�:�;�8�e�L���YӖ��V��C1��*���d�l�
�a�k�}��������l0��h��D��
�f�d�u�8�3���B�����R�����!�<�3�
�`��E��Yے��lR��E��G��u�:�u�%�4�3����H���9F������!�&�3�
�f��E��Yۋ��l0��B1�B���u�;�u�8��i����H¹��]ǻN��*���g�d�
� �����Lù��Z�=N��U���u�%�6�;�#�1�Fف�?����[�������
�
�
�
�"�l�Eف�K���F�G�����_�u�u�u�w�����Mǹ��l_��h����u�
�4�g�f��(�������G9��h_�M���u�h�_�u�w�}�W�������l
��h^�����}�8�
�
�d�/���L����[�I�����u�u�u�u�w�<�(���
����9��=N��U���4�g�d�
�"��(���H����CU�
NךU���u�u�%�6�9�)���&Ġ����YN�����2�
�
�d�>�;�(��M����O�I�\ʰ�&�u�u�u�w�}��������l ��^�*��_�u�u�
�6�o�F�������
P��N�U���u�u�u�4��2�����Г�V��@��U �1�'�9�"�f�;�(��A����O�I�\ʰ�&�u�u�u�w�}��������l ��^�*��_�u�u�
�6�o�Eہ�&����l��C1��*��m�%�u�h�]�}�W���Y����\��h��*���=�;�}�8��l�Eہ�����V�N��R��u�9�0�_�w�}�W���	����@��A[��N���u�%��9�����L����[�N��U���!�%�g�
�"�n�N���Y����N��G1�����c�
�g�e�w�}�F�������9F�N��U���
� �a�f�'�f�W���	����9��h��G���%�u�h�'��;�(��&����F�G1��؊�d�3�
�f��l�K���)����U��Z��D��x�d�1�"�#�}�^�ԜY�Ƽ�e��h]�����f�
�g�i�w�)�(�������P������� �&�2�0��)�(�������P�������%��9�
�f�;�(��&���F��P ��]��u�%��9��l����JĹ��O�\�\�ߊu�u�
�4�e�n�(���O�ߓ�F������f�
� �g�`�-�_������\F��d��Uʥ��9�
�a�1��Bށ�K���@��[�����6�:�}�;�>�3�Ǯ�/���� U��B1�L���|�~� �&�0�8�_���&�ӓ�l �� Z�����n�u�u�%��1�(�������9��R�����g�3�
�m��o�}���Y����_T��1��*��
�d�i�u���(���O�ғ�N��N����!�u�|�_�w�}�(���K����U��_��G��u�!�
�:�>�����۔��Z��B �����}�!�
�:�>�����ە��]��G1��؊�m�3�
�a��m�W�������A��H��#���
�m�3�
�c��F���U����]ǻN��*���g�f�3�
�g��E��Y����_	��T1�����}�;�<�;�3�-�!���&����T9��[��^ʠ�&�2�0�}�:��F���&����CW�d��Uʥ��9�
�e�1��A݁�M���C9��[\��M���
�a�
�g�e�}�������9F������a�
� �m�c�-�W��
����\��h����� �&�2�0������Mù��lQ��h�U���;�<�;�1�#�-�E߁�&����V��G����u�
�4�g�c����@����[��C
�����
�0�!�'�"�.����Q����_T��1����l�|�~� �$�:��������l��B1�C���|�n�u�u�'��݁�N����V��h�I���!�
�:�<��8��������]��G1��؊�c�'�2�g�f�t�\ϫ�
����WN��G1�*��� �d�b�
�f�t�}���Y����_T��h��D��
�f�i�u�w�}�W���	����9��h��D��
�f�"�0�w�)���&����lW��1��]���h�r�r�u�;�8�}���Y���A9��\�� ��b�
�d�_�w�}�(���K����U��Z�����h�_�u�u�w�}�(�������9��h_�E���u�=�;�}�:��(������� S��G��U��|�0�&�u�w�}�W�������9��h_�A���n�u�u�%��1�(�������
T��N�U���u�u�u�%��1�(�������G9��D�� ��f�
�f�"�2�}����L¹��U��X�����|�h�r�r�w�1��ԜY���F��e�����`�3�
�f�e�-�L���YӖ��R
��]�� ��a�
�f�i�w�}�W���YӖ��R
��\�� ��l�
�f�"�2�}����L����U��_�����|�h�r�r�w�1��ԜY���F��e�����c�3�
�a�o�-�L���YӖ��R
��[�� ��e�
�f�i�w�}�W���YӔ��lW��Q��A���%�u�=�;��0�(�������R��F�U���d�|�0�&�w�}�W���YӖ��R
��1��*��c�%�n�u�w�-�!���&ƹ��lW��1��U��_�u�u�u�w�����M����R��h����u�!�%�`�����H˹��V�
N��R���9�0�_�u�w�}�W���&�Փ�F9��Z��D�ߊu�u�
�4�e�k�(���H����CU�
NךU���u�u�
�0�"�)�D݁�����9�������8�
�d�g��8�(��I���F�G�����_�u�u�u�w��(�������R��UךU���
�4�g�c��(�F��&���FǻN��U���
�4�g�g����������U��Y�����=�;�}�8��o����&����l��G��U��|�0�&�u�w�}�W���	����F
��]�� ��g�
�a�_�w�}�(���K����U�� V�����h�_�u�u�w�}�(���K����U�� ]�����=�;�}�8��n����&����l��G��U��|�0�&�u�w�}�W���	����F
��Z�� ��b�
�a�_�w�}�(���K����U��Z�����h�_�u�u�w�}�(���A����^��h����u�!�%�b��(�F��&���F�_��U���0�_�u�u�w�}�(���K�ѓ�F9��X��F�ߊu�u�
�4�e�k����N�֓� F�d��U���u�%��9��l����O�ӓ� F��R �����c�
�
� �f�m�(��I���W����ߊu�u�u�u���A���&����l��=N��U���4�g�b�3��j�A���Y���F�N�����9�
�
� �f�i�(��������hX�����
�b�m�%��t�J���^�Ʃ�@�N��U���'��d�
�"�l�@ہ�H���F��a��*��� �d�`�
�d�a�W���Y�����T�����d�
�e�e� �8�Wǫ�����\��B1�Gڊ�g�e�u�u�f�t����Y���F������a�
� �l�n�-�L���YӖ��9��h\�C���u�h�}�
�b�j�E���&����R����U���7�'�'� �3�+��������l ��_�*��n�u�u�%�>�;�(��K����[�G1�B݊�
�
�0�
�d�j��������A9��B �����9�"��3��m�N���P���F��Y��ۊ�
� �d�g��o�K���
����Z��h��*��l�-�'�6�%�$�F���&����l��d��Uʥ�;�!�<�<�1��Nށ�K�����Y��*���
�g�`�-�%�>��������9��UךU���
�%�3�
�o��E��Y����_	��T1�����}�;�<�;�3�)���&����U��G��U���<�;�1�4��2����Ź��]ǻN��*��� �a�f�%�w�`�}���Y���R��X ��*���c���u�?�3�_�������lT��h�E���u�d�|�0�$�}�W���Y����C9��Y����
�n�u�u�&������ד�F9��1��U��}�
�
�
�"�h�B���Y����B��R	��G��n�u�u�$��.����J����R��G\��H���
�
�
�
�"�j�B���Y����B��h��B���%�|�_�u�w�?��������U��Z��G��u�'�<�<�����A����R��F��*ۊ� �b�g�%�~�W�W�������Z�� 1��*��
�g�i�u�#�-�C؁�����l��V �����
�
� �m�e�-�^�ԜY�ƽ�l��^	��L���
�f�
�g�k�}����L����l_��h����$�<�
�
�"�d�G���P���F��h��A���%�u�h�_�w�}�W���
����U��]��Fʢ�0�u�!�%�f����J����O�I�\ʰ�&�u�u�u�w�}����Kʹ��lR��h����u�7�!�d�1��@݁�J���C9��[\��M���
�a�
�g�b�9� ���Y����F�F��*؊� �m�g�%�w�`����J����T��G\��U���u�:�;�:�g�f�W������� 9��hW�*��i�u�
�
�g�;�(��&���K�
�����e�n�u�u�&�4�(���N�ߓ� F������f�
� �g�`�-�_�������S�=N��U���
� �b�d�'�}�J���[ӑ��]F��Z��L���
�d�
�d�j�<�(���
����9�������w�_�u�u�����M����[�L�����}�8�
�g�1��O߁�H����C9��Y�����e�u�9�0�u��}���Y����V��B1�C���u�h�&�1�;�:��������@��R
�����l�<�3�
�o��F���Y����V��Z��B���3�
�b�
�f�t�}���Y����W��B1�Fފ�d�i�u�!��2����������^�� ���2�0�}�
�����KĹ��J��G�U���'��d�
�"�l�@ׁ�H���@��[�����6�:�}�0�>�8��������A9��1��*��m�%�|�a�~�f�W������� 9��h_�A���u�h�&�1�;�:��������A��M�����;�1�'��a�;�(��M����R��UךU���
�
�a�3��i�E���Y����G��X	��*���!�'�'�&�-�u��������l0��h��D��
�a�y�e�~�W�W���&����l ��X�*��i�u�!�
�8�4�(�������V��RF�����0�}�
�
��(�F��&���V�d��Uʧ��d�
� �f�l�(��E�ƿ�W9��P�����:�}�0�<�2�(�����ξ�e9��Q��B���%�|�a�|�l�}�WϬ�/����U�� Y�����h�&�1�9�0�>�����ξ�@�������1�'��&�1��@���	���O�=N��U���
�m�3�
�o�o����Dӕ��l
��^�����'�'�&�/��3����۔��lW��B1�D؊�a�y�e�|�]�}�W���&¹��lW��1��U��%��9�
��(�F��&���
F��@ ��U���_�u�u�
�����J����[��C
�����
�0�!�'�$�:��������l��B1�@���|�x�&�2�2�u����J����F9��1��\��u�u�'��d�;�(��&���F��S1�����#�6�:�}�>�3�Ǫ�	����Z9��hV�*��u�u�<�;�3�)���&����l^��h�\�ߊu�u�
�
��(�F��&���F��B�����&��'�2�e�i�W���	����@��A_��E��u�u�'��b�;�(��A����[��h8��G���
� �d�a��n�D�������R�=N��U���
�
� �d�e��C��Y����_T��h��D��
�f�f�u�8�3���B�����hY�� ��b�
�a�i�w�����L����R��h�F���:�;�:�d�l�}�WϬ�/�ޓ�F9��Y��F��u�;�8�0��?�(���&����U��H�����;�!�9�d��t�}���Y����
9��h_�M���u�h�%��;��F���&����l��W�����:�a�n�u�w�/�!���&����CT�
N�����2�6�#�6�8�u����ے��lW��^1��*��
�d�u�u�>�3�Ǫ�	����Z9��hX�*��|�_�u�u���(���H����CR�
N��#���
�
� �d�c��D��Y����G	�UךU���
� �`�l�'�}�J�������l ��X�����;�u�8�
�n�;�(��&���9F���*���<�3�
�l��o�K������� 9��hY�*��:�u�
�
�"�j�C���P���F��^1�����l�
�g�i�w�)���&����T�������2�g�f�|�]�}�W���&����U��[��G��u�!�%�a��(�@���	�ƣ���h��B���%�|�_�u�w�8�(���Hù��l ��W�*��i�u�&�9�#�-�(�������^��N��ʻ�!�&�9�!�'��F���&����l��d��Uʦ�9�!�%�e�>�;�(��K����[�D�����
�
� �d�g��DϿ�ӈ��l��h��L���3�
�c�c�'�t�}���Y����G��1�����4�
� �`�`�-�W��Q����G��h
�����;�3�
�`��o��������F9�� 1��\�ߊu�u�0�
�:�l�(�������^��N�U¦�9�!�%�
�f�;�(��M����R��C��C܊�d�3�
�m�o�-�^�ԜY�ƿ�_9��G_�����
�c�m�%�w�`�_���&����l��B1�Mފ�g�4�1�!�'�h�(�������9��UךU���0�
�8�d�1��Dց�K�����h_�� ��`�%�u�:�w�-��������lW�=N��U���
�8�d�<��(�F��&���F��Z��A���3�
�m�g�'�}����	����@��A_��\�ߊu�u�0�
�:�l����&����l��S�����`�
�
� �f�l�(������C9��Y�����d�n�u�u�$�1����&����S��N�U¡�%�`�3�
�b��EϿ�ӕ��l��1��*��
�g�n�u�w�.����	����l ��W�*��i�u�!�%�a��(���H����CT��Y
�����8�d�<�
�"�l�Fׁ�K��ƹF��R�����<�3�
�`�c�-�W��Q����R��h��D��
�g�4�1�$�1����&����lW��1��\�ߊu�u�0�
�:�n����L¹��Z�=N��U���u�8�
�a�1��A܁�Hӑ��]F��R�����3�
�a�
�e�m�W���H����_��=N��U���u�%�6�;�#�1�Fف�B�����h��F���
� �d�f��o�K�������9��h��D��
�g�-�'�6�����&����O��N�����!�%�
�
�"�l�N߁�K�����h[�����
�`�m�%�w�2�W�������l
��h_����u�0�
�8�c�;�(��&���F��T��*���f�f�%�u�9�}��������lS��h�N���u�&�9�!�'��F���&����l��S�����c�3�
�l�a�-�W���Y����G��h�����l�a�%�|�]�}�W���&����l��B1�E؊�g�i�u�!�'����@Ź������*���g�<�3�
�b�i����s���@��C��*���:�2�;�3��h�(��E����^��h��F���%�u�'�!�'�h����LĹ��]ǻN�����8�c�3�
�a��E��Yە��l��1�����4�
� �`�n�-�W���Y����\��h��*���_�u�u�0��0�A���&����
R��G]��H�ߊu�u�u�u�:��N�������Q��N�����&�9�!�%��l����@�ԓ�N��S��D���0�&�u�u�w�}�Wϭ�����l��Q��L���%�n�u�u�$�1����&����lW��1��U��_�u�u�u�w�0�(�������S��h����u�&�9�!�'��(���H����CT�N��R��u�9�0�_�w�}�W�������C9��Q��@���%�n�u�u�$�1����&����W��N�U¼�8�
� �f�`�-�W���Y����G��h��@���%�|�_�u�w�8�(���A����W��G]��H�ߊu�u�u�u��<�E�������9�������0�
�8�b�%�:�E��Q���A��N�����u�u�u�u�$�1����&����T��d��Uʦ�9�!�%�3��e�(��E����V
��Z�*���:�2�;�3��j�(������C9��Y�����d�n�u�u�$�1����¹��lW��1��U��}�8�
�a�>�;�(��K����R��Y�����0�1�:�;�2��(ށ�����P�=N��U���
�8�
�
�"�l�@܁�K�����h[�����
�`�g�%�w�3�W�������V��X�����
�0�
�f�`�f�W���Y����[9��C1����� �f�f�%�w�`��������l��C�����/�}�<�;�3�.�(���&����S��G�G���_�u�u�&��0�(���J�ӓ� F�d��U���u�!�%�f�1��D܁�Kӑ��]F��T�����g�
�g�e�w�}�F�������9F�N��U���
�
� �f�n�-�L���Yӕ��T
��G�����;�3�:�!�2�-�!���H����W��h�I���!�
�:�<��8��������]��C��Bۊ�
� �g�a��l�W�������V��G1�����9�m�b�|�l�}�Wϭ�����C��^�����:�!�0�%��4����I�ד�F���*���<�
�0�!�%�(�����θ�C9��h�� ��f�
�d�u�w�3����ۇ��P	��C1��M��|�n�u�u�#�-�(���H����CT�
N�����9�"�3�
�g�o����ӈ��l��h ��*��� �d�f�
�e�f�W�������l ��W�*��i�u�!�%�a��(���H����CT��Y
�����8�f�<�
�"�l�D߁�K��ƹF��Z�����d�c�%�u�j�u��������l ��_�*��:�u�0�
�%��(���&����lW��1��\�ߊu�u�8�f�1��B���	���N��G1�*��� �d�f�
�e�<�ϭ����� 9��Q��@���%�|�_�u�w�}�W���&�֓�F9��1��U��&�1�9�2�4�+����Q����I��^	��¡�%�d�
� �d�n����J���9l�N��Uʡ�%�d�
�
�"�k�F���Y����G��X	��*���!�'�'�&�-�u����ۍ��A9��F_��D���n�_�u�u�:��F���&����CR�
N��*���f�d�%�}�f�9� ���Y����F�N�����d�
�
� �a�h����Dӕ��l
��^�����'�'�&�/��4��������9��B�\��_�u�u�8��o����Hƹ��Z�D�����6�#�6�:��5��������]��Y�����d�
� �a�f�-�^ê�&����T��B �����}�e�u�u�?�<����
����lU��h�F���u�:�;�:�g�t�^��Y���F��Z��G���3�
�b�
�f�a�W���&����P9��T��]���<�0�&�2�2�u����K����W��UװU���!�%�d�
�"�i�D���Y���D��_��]���;�1�!�%�d�;�(��&���F��P ��]���6�;�!�9�f��A�������V�=N��U���u�8�
�f�>�;�(��&���F��S1�����#�6�:�}�2�4�ǭ�����X��h\��E���b�|�_�u�w�)���&����U��N�U���
�
� �g�`�-�_��T����\��XN�N���u�!�%�d��(�C���	�����h�����0�!�'� �$�:����K���� W��G\��^ʠ�&�2�0�}�'�>��������u ��UךU���8�
�`�<�1��C؁�H���@��[�����6�:�}�0�>�8��������B��D�����3�
�a�
�e�q�@���s���G��X�� ��`�%�u�h�u�� ���Yە��]��q\�� ��d�%�|�k�$�:����	����@��A_��D���u�9�0�w�u�W�W�������l ��Y�����h�&�1�9�0�>�����ι�@��R
��G���
�d�
�g�w�}��������C9��Y����
��|�n�w�}����H˹��lR��h�I���d�u�=�;��4��������9��hZ�*��u�u�<�;�3�<�(���
����T��G�����u�e�n�u�w�)���&����U��N�U��u�=�;�}��8����
����W��G\��U���6�;�!�9�b��^ϻ�
���]ǻN�����
� �f�`�'�}�J���[ӑ��]F��Z��*���g�l�%�u�w�-�������� 9�������w�_�u�u�:��G���&����CR�
N��*���
� �f�`�'�u�FϺ�����O��N�����g�
�
� �o�m����Dӕ��l
��^�����'�'�&�/��3����ۗ��R��P ��*���m�a�%�|�f�t�L���YӒ��lT��Q��Eފ�d�i�u�!��2����������^�� ���2�0�}�7�6�.����&����
_��G�C���_�u�u�8��n����@ʹ��Z�C��C���
�l�
�g�f�}�W�������V�=N��U���
�a�3�
�g�e����D���F�N����
� �g�`��l� ���Yۖ��Q��1�����g�l�}�|�j�z�P������F�N�����g�
�0�
�c�d�}���Y���G��Z��*���m�e�%�u�j�.��������V��EF�����}�<�;�1�<�/�(ށ�I����O��=N��U���u�8�
�`�>�;�(��&���F��S1�����#�6�:�}�2�4�ǭ�����C9��[\��A���
�`�
�g�{�e�^�ԶY����^��1��*��
�d�i�u�:��E���&����CT�N�Dʱ�"�!�u�|�]�}�W���&�ѓ�F9��\��F��u�u�u�u�w�)���&����S��G_�����}�
�`�b�e�4�(���&����V�
N��R���9�0�_�u�w�}�W���&�ӓ�V��]����u�8�
�m�>�;�(��&���F��S1�����#�6�:�}�2�4�ǫ�
����WN��h�����b�'�2�g�g�t�F���B�����h\�����a�
�f�i�w�<�(�������l��C�����0�}�;�<�9�9����@¹��@��B1�@���|�u�:�;�8�)�(�������F��P ��]���
�d�6�&��(�C���	�����YN�����!�2�'� �$�:��������l��C1��*��
�d�|�h�g�<�Ϫ�&����T��B �����}�8�
�d�4�.�(���M�ӓ�O�
[�U���0�w�w�_�w�}����&����_��N�U���2��3�
�c��F��Y����W	��C��\�ߊu�u�8�
�����J����[��C
�����
�0�!�'�%�.��������V��Z��C���3�
�g�
�c�q�C���s���G��^�� ��f�%�u�h�#�-�F؁�����l��N�Dʱ�"�!�u�|�]�}�W���&�ד�F9��1��U��_�u�u�u�w�-��������lU��@��U¡�%�d�
� �c�j����P���A�R��U���u�u�u�%�8����N����9F���*���3�
�e�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���&�ד�F9��1��\���|�n�u�u�#�-�D݁�&����T��N�U»�"�<�;�<��(�N���	�ƴ�AF��h�����#�
�|�_�w�}����J����V��G\��Hʦ�1�9�2�6�!�>��������_�������1�4�
�:�$�����J����u ��q(��3���:�<�!�2�%�(�������F�C��F؊� �`�d�%��l�FϺ�����O�G�U���!�%�f�
�"�h�F���Y���G��]�� ���`�%�u�:�w�-��������9��q(��3�����|�_�w�}����M����F9��1��U��}�<�;�<��8�(��LӞ����T�����d�d�n�u�w�)���&���� S��N�U���4�g�g�3��o�(��H�����Y��E��u�u�!�%�d��(���@�֓�F�F�����;�<�
� �n�i����Ӗ��V��C1�����3�
�b�
�e�f�W�������9��hX�*��i�u�-�
�2�0�(���?����c	��C1��#���
�d�
�f�a�p�FϺ�����O��N��U���!�%�f�
��(�O���	�����h�����0�!�'�'�$�'�_�������R��1��\��|�n�_�u�w�0�(�������9��R�����9�
�d�3��n�(��L�����Y��E��u�u�u�u�#�-�Dց�&����T��N�U���
�:�<�
�2�)�Ǭ�
����@��R
��*���g�a�
� �o�i����H���9l�N�����3�
�f�
�e�a�W���&����P9��T��]���<�;�1���(�D���	�����^	��´�
�:�&�
�!�o�1��P���F��G1�*���b�b�%�u�j�-�!���&�ד�F9�� 1��]���:�;�:�c�l�}�WϪ�	����U��^��D��u�
�4�g�d����H����F�N�����u�|�_�u�w�0�(�������V��h�I���!�
�:�<��8��������VN��D�����7�4�&�2������J���P�d��Uʡ�%�a�
� �`�m����DӖ��R
��V�� ��d�%�}�u�8�3���B�����hZ�����
�e�e�%�w�`�_���
����Z��h��D��
�f�-�'�6�����&����O��N�����a�
� �m�c�-�W������l ��\�����u�:�;�:�f�f�W�������9��Q��D���%�u�h�}�>�3����&����U����U���6�;�!�9�f�l�L���YӒ��lR��B1�L���u�h�&�1�;�:��������F��P ��]���6�;�!�9�f��^������]��q\�� ��d�%�|�n�w�}����Lù��U��_�����h�}�0�&�0�?��������T��N��U���0� �!�c�9�)����&����l��d��Uʡ�%�`�
�
�"�l�A݁�K���W�@��U¥��&�9�
�c�4����J�ԓ�F�V�����
�#�
�|�2�.�W��B�����h[�����g�
�f�i�w��(�������9��_�����:�d�n�u�w�)���&����lW��1��U��w�w�"�0�w�-�%�������l��B1�EҊ�a�h�4�
�8�.�(���&����_��^�����u�8�
�f�>�;�(��K����[�L�����}�
�`�d�d�4����M�Г� F�V�����
�#�
�m�w�1����[���F��G1�*���d�d�
�f�k�}��������V��_��#���
�e�c�%��h��������]ǻN�����a�<�3�
�b�e����D������YN�����;�1�%�e�o��(�������9��N� ���2�0�}�%�4�3����L����F��D��E��u�u�!�%�b��(���H����CT�
N��Wʢ�0�u�;�8�2�� �������_$��D1�����`�a�%�u�w�-��������lU�R��U��n�u�u�!�'�h�(�������9��R��W���"�0�u�;�:�8�(���:����P��^��#���
�`�a�%�w�}��������ET��N�����e�n�u�u�#�-�B؁�����9��R�����9�
�
� �f�h�(��K�ƨ�D��\�N���u�!�%�`�����OĹ��Z�^�����u�%��&�;��O���&����l��
N��*���&�
�#�c�g�}����[����F�C��@ӊ� �d�`�
�f�a�W�������Q��h��D��
�f�g�x�f�9� ���Y����F�C��@ӊ�
� �g�d��l�K�������T��A�����0�<�0� �$�:��������l��Y
�����:�
�
� �e�m�(��U���9F���*ߊ� �f�b�%�w�`�U������� ��Q��Dۊ�g�h�4�
�8�.�(���K���V
��L�N���u�!�%�c�����JĹ��Z�D�����6�#�6�:��8��������]��G1�Mۊ�
�
� �g�e��D��P��ƹF��Z��D���
�`�e�%�w�`��������l��C�� ���2�0�}�
�b�l�D�������
P��G��U���<�;�1�4��2����ƹ��]ǻN�����d�<�3�
�g�n����DӖ��V��C1�*���g�m�
�`�]�}�W���&�ԓ�F9��X��D��u�!�
�:�>�����۔��Z��B �����}�8�
�d�1��B���	���O�=N��U���
�g�<�3��j�E���Y���D��_��]���0� �!�g�����@����[��G1�����9�a�e�u�;�8�U���s���G��]�� ��`�
�g�i�w�)�(�������P�������0�!� �&�0�8�_�������l
��1��3���!�
�;�0�2�u�������A���*���3�
�`�c�'�u�A������\F��G��N���u�!�%�c�����L˹��Z�_�����u�%��&�;��@�������^��N�����:�&�
�#��t����Y���9F���*���3�
�`�c�'�}�J�������l ��[�*��-�'�4�
�8�.�(���O����uO��N�����c�
�
� �f�h�(��E���F��R ����m�
�
�d�1��O���	���R��X ��*���
�m�u�9�2��U�ԜY�Ƹ�C9��h�� ��`�
�g�i�w�l�W����ι�@��R
��*���d�f�<�
�"�l�Dف�J���F��P ��]���6�;�!�9�b�l�^������D��N�����c�
�d�3��e�O���Y���D��_��]���7�'�!�:�%�)��������lW��B1�Cފ�d�h�4�
�8�.�(���&����_��^�����u�8�
�c�>�;�(��&���F��G1������
�<�0��4����/����W��G]��@ʱ�"�!�u�|�]�}�W���&�ѓ�F9��Z��D��u� �7�'�%�(��������lR��B1�Eي�g�g�u�u�w�2����I��ƹF��Z��B���3�
�m�a�'�}�J���[ӑ��]F��B�����:�'�!�6�;�4����H����^��h�Hʴ�
�:�&�
�!��^ϻ�
���]ǻN�����m�3�
�g�e�-�W������\��C��*��
�
� �d�g��D��Y����G	�G�U���!�%�c�
��(�F��&���F�N�����%��&�9��k����@�ԓ�F�V�����
�#�c�e�w�1����[���F��G1�����l�
�g�i�w�)�(�������P�������<�=�}�<�9�9����/����_��G]�����;�0�0�}�9�4����^�����hW�� ��l�%�}�d�f�9� ���Y���O��N�����c�<�3�
�b��F��Y����_	��T1�����}�0�<�0�"�.����Q����}"��v<�����d�
� �c�n�-�^��P��ƹF��Z��E���3�
�d�d�'�}�Jϭ�����Z��R��§�&�/�}�;�>�3�ǰ�����A	��S!�����"��d�3��l�D���P���l�N����
� �d�e��n�K���&����lQ��B1�L܊�f�g�u�:�9�2�E���s���G�� _��*���g�a�
�d�k�}��������E��X�����0� �&�2�2�u�(��H�ғ�9��h\�E���|�m�|�_�w�}����K����F9��Y��D��u�
�0� �#�n�(���K����CS��N�����b�
� �d�f��F��Y����V��U��*ߊ� �d�m�
�d�o�Z������\F��d��Uʡ�%�b�
� �f�e�(��E�ƿ�W9��P�����:�}�;�<�9�9���A¹��ZW��B1�F܊�f�u�u�;�>�3�ǿ�&����G9��1�\�ߊu�u�8�
�a�;�(��O����[��C
�����
�0�!�'�%�.��������V��Z��@���
�m�e�%�~�l�^��Y����^�� 1��*��e�%�u�h�$�9��������G	��D�����3�}�;�<�9�9��������_��h(��3���:�<�!�2�%�(�������F�C��B܊� �d�m�
�f�l�Z�������V�G����u�8�
�m�1��O���	���N��G1�*���d�l�
�g�/�/��������_��h(��3��u�u�!�%�`�;�(��&���F�N����� �&�2�0��5��������9��N� ���2�0�}�%�4�3����H����O��[��W���_�u�u�8��l����H�ޓ�F� �����'� �1�0�"�)�!�������Q��F�U���u�:�;�:�g�f�W�������l ��Y�����h�<�0�
��(�E���	����K�
�����e�n�u�u�w�}����@¹��@��B1�@���u�h�&�1�;�:��������A��M�����1�!�%�d��(�C���	���O�=d��Uʡ�%�l�3�
�o��F��Y����_	��T1�����}�0�<�0�"�.����Q����^��V�����`�
�d�y�c�t�}���Y����U�� W��F��u�4�
�:�$��ށ�Y�Ƹ�C9��Q��Bߊ�d�n�u�u�#�-�ށ�M����U��h�I���d�u�=�;����������U��W�����u�%�6�;�#�1�O��Y����D��d��Uʡ�%�<�
� �f�k�(��E���F��R �����;�1�
�0�:�l�B�������R��N�����:�&�
�#�a�m�W�������l�N�����g�
� �d�b��E��Y���D��F��'���9�
�d�3��o�G���Y�ƭ�l��D��Ҋ�|�0�&�u�g�f�W�������l ��\�*��i�u�d�u�?�3�_���&����l��Z1�L���3�
�e�c�'�}�W�������l
��1�U���0�w�w�_�w�}����&����W��N�U���
�:�<�
�2�)�Ǭ�
����F��P ��]���
�8�
�
�"�o�F���P����]ǻN�����3�:�
�
�"�l�Bׁ�K�����h��*ۊ� �d�g�
�e�<�ϼ�����V��1�����d�g�%�|�]�}�W�������D9��h_�E���u�h�}�0��/�(���@�Г�F��SN�����0�e�<�<�1��G���	����V��U����