-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�u� �2�4��������T��_�[���n�_�&�u�2�8��������l��^	��Ĵ�9�_�0�!�#�}�1��@����lV��hW�����c�'�8�<�w�}�WϹ�����l�N��U���u�u�"�1�?�}�W������V�
N�N�ߊu�u�u�u�w�}�������F��^ �����o�u�f�u�w�}�W���Y���^��D��U���o�<�!�2�%�g�W��N���O��=N��U���!�}�u�u�w�}�WϿ����F�N��U���
�:�<�
�2�)�ǿ�����F��@ ��U���u�u�u�u�w�}���Y���\��YN�����2�6�u�u�w�}�W������F�N����&�1�9�2�4�+����Q����G�
�����e�n�u�u�w�}�WϽ����F������9�2�6�u�w�t�W��Ӄ��Z��dװ���<�0�!�'�w�)�W�������
'��Q1�����>�'�
�
�8�}��Զ
����_F��S�����o�&�1�9�0�>�����έ�Z��_�����:�e�n�_�.�8����������V�����u�:�8�8�$�'�Z����ƿ�W9��P�����:�u�1�<�#�p�W������]�D�����0�u�u�0��/����D��ƹF�S�W��e�e�e�e�g�m�G��I����V��^�W���u�u�d�h�w�m�F��I����W��^�E��d�d�d�e�g�q�}���Y���D��_�D��e�d�e�e�g�l�F��I����D�=N��U���k�w�e�d�g�m�G��H����V��_�D��d�w�u�u�w�i�J���I����W��^�E��e�e�d�d�f�l�F��U���F��
P��E��d�d�d�d�f�l�G��I����V��_�Y�ߊu�u�u�k�u�m�F��H����W��_�D��d�e�d�d�u�}�W���N���V��_�D��e�d�d�d�g�l�F��H����J�N��M��u�e�d�d�f�m�G��I����W��_�E��e�y�_�u�w�}�I���I����W��^�D��d�e�e�d�f�l�G���Y���W��
P��E��d�d�e�d�f�l�G��I����W��^�Y�ߊu�u�d�h�w�m�F��H����W��^�D��e�d�e�e�f�q�}���Y���F�_�E��e�d�d�e�f�m�G��H����W�d��U��u�k�w�e�f�m�F��I����W��_�D��e�e�w�u�w�}�F���G����W��_�D��d�d�d�d�g�l�F��I���9F�_�H���e�d�d�d�f�l�F��I����W��^�E��y�_�u�u�a�`�W��H����W��_�D��e�d�d�e�g�m�G��s���Q�	N��E��e�d�d�d�f�l�G��I����W��_��U���u�d�u�k�u�m�F��H����V��^�E��e�d�e�e�u�}�W���H���D��_�D��d�d�d�d�g�m�F��I����D�=N��U��h�u�e�d�f�l�F��H����V��_�E��e�e�y�_�w�}�F��Y����W��^�E��d�d�d�e�g�m�G��I���F�\��K���e�d�d�e�g�m�G��I����V��_�D���u�u�u�g�w�c�U��H����V��^�D��e�d�d�d�f�l�U���Y���F�L�D��e�e�e�e�f�l�G��H����W��L����u�`�h�u�g�l�F��I����V��^�E��d�e�d�d�{�W�W���O���V��_�E��e�e�d�d�f�l�G��H����J�N��G���k�w�e�d�f�m�G��I����V��^�E��d�w�u�u�w�o�W���[����W��^�D��d�d�d�e�g�m�G��[��ƹF�N��U��d�d�e�e�f�m�F��H����V��_�E���_�u�u�e�j�}�G��H����W��^�D��d�d�d�e�f�m�[�ԜY����[�^�D��e�d�e�e�g�l�G��I����W��B��U���f�u�k�w�g�l�F��H����W��^�D��e�e�e�w�w�}�W��Y���V��_�E��d�d�e�e�g�l�F��H����FǻN��A��u�e�d�d�g�m�G��I����W��^�E��e�y�_�u�w�h�J���I����V��^�E��d�e�d�d�g�m�F��U���F��S�W��d�d�e�d�g�m�G��I����W��_�W���u�u�f�u�i��G��H����V��^�D��e�e�e�e�f��W���Y����X�^�D��e�d�d�d�f�m�G��H����W��NךU���l�h�u�e�f�l�G��H����V��_�E��d�d�e�y�]�}�W��D���W��^�D��e�d�d�d�g�l�F��I���l�N�U��w�e�d�d�g�m�G��I����W��_�D��w�u�u�u�c�}�I���I����V��^�D��d�e�e�d�f�m�F���Y���R��
P��E��d�e�d�e�g�l�G��I����V��_�Y�ߊu�u�a�h�w�m�F��I����W��^�D��d�e�d�e�g�q�}���Y���F�_�D��e�e�d�d�f�l�F��H����V�d��U��u�k�w�e�f�l�G��H����V��^�E��d�d�w�u�w�}�C���G����W��^�E��d�d�d�e�g�l�G��I���9F�Z�H���e�d�d�e�f�m�G��H����V��_�D��y�_�u�u�n�`�W��H����W��_�D��e�d�d�d�f�m�G��s���V�	N��E��d�e�e�d�f�l�G��I����V��^��U���u�`�u�k�u�m�F��I����V��^�E��e�e�e�e�u�}�W���L���D��_�E��d�e�d�e�g�l�F��I����D�=N��U��h�u�e�d�f�m�F��I����W��_�E��e�e�y�_�w�}�C��Y����W��_�E��d�e�e�e�g�l�G��I���F�[��K���e�d�d�e�g�m�F��H����V��_�E���u�u�u�`�w�c�U��H����V��_�D��d�d�e�d�f�m�U���Y���F�L�D��e�d�d�e�f�m�G��H����W��L����u�m�h�u�g�l�F��H����W��_�E��e�e�d�e�{�W�W���@���V��_�E��d�e�d�d�f�l�G��H����J�N��C���k�w�e�d�f�m�G��H����W��^�E��d�w�u�u�w�k�W���[����W��^�D��d�e�d�d�f�l�G��[��ƹF�N��U��d�d�e�d�g�m�F��I����W��_�D���_�u�u�f�j�}�G��H����V��^�D��d�e�e�e�f�l�[�ԜY����[�^�D��e�d�e�e�f�m�G��I����V��B��U���c�u�k�w�g�l�F��H����V��^�D��d�e�e�w�w�}�W��Y���V��_�D��d�d�e�e�g�l�F��H����FǻN��B��u�e�d�d�g�l�G��H����V��_�E��d�y�_�u�w�e�J���I����V��^�D��e�d�e�e�g�m�F��U���F��S�W��d�d�e�d�f�m�G��H����V��_�W���u�u�b�u�i��G��H����W��_�D��d�d�e�e�g��W���Y����X�^�D��d�e�d�d�g�m�G��H����V��NךU���g�h�u�e�f�l�G��H����V��_�E��d�e�e�y�]�}�W��D���W��^�D��d�d�d�e�f�m�F��I���l�N�U��w�e�d�d�g�l�G��I����V��_�D��w�u�u�u�`�}�I���I����V��^�D��e�e�d�e�g�m�F���Y���Q��
P��E��d�e�d�d�f�l�F��H����W��^�Y�ߊu�u�b�h�w�m�F��I����V��_�D��e�e�d�e�f�q�}���Y���F�_�D��d�d�d�d�g�m�G��H����V�d��U��u�k�w�e�f�l�G��H����V��_�D��d�d�w�u�w�}�O���G����W��^�D��d�e�e�d�g�l�F��H���9F�V�H���e�d�d�e�f�l�F��I����V��^�D��y�_�u�u�e�`�W��H����V��^�E��e�e�e�e�f�m�F��s���U�	N��E��d�d�e�e�g�m�F��I����V��_��U���u�m�u�k�u�m�F��H����V��_�D��d�e�e�e�u�}�W���A���D��_�E��e�e�e�e�f�l�F��H����D�=N��U��h�u�e�d�f�m�G��I����V��^�D��e�e�y�_�w�}�@��Y����W��^�E��e�e�e�e�g�l�G��H���F�V��K���e�d�d�d�g�m�G��I����V��^�D���u�u�u�m�w�c�U��H����V��^�D��e�d�e�e�g�l�U���Y���F�L�D��e�e�e�d�g�m�G��H����V��L����u�d�h�u�g�l�F��I����W��_�E��d�d�e�e�{�W�W���K���V��_�D��d�e�e�d�f�m�F��H����J�N��L���k�w�e�d�f�l�G��I����V��_�E��d�w�u�u�w�d�W���[����W��^�E��d�e�d�d�g�l�G��[��ƹF�N��U��d�d�e�e�g�m�G��H����V��^�D���_�u�u�c�j�}�G��H����V��_�D��e�d�e�e�f�m�[�ԜY����[�^�D��d�e�d�e�g�l�F��H����W��B��U���l�u�k�w�g�l�F��I����W��^�D��e�d�e�w�w�}�W��Y���V��_�E��d�d�e�d�f�m�F��I����FǻN��E���k�w�e�d�f�l�G��H����V��^�E��e�w�u�u�w�l�F��Y����W��^�D��e�e�d�d�g�l�F��H���F�^�H���e�d�d�e�g�l�G��I����W��_�D��y�_�u�u�g�}�I���I����W��^�E��d�d�d�d�f�l�G���Y���W��S�W��d�d�d�e�g�m�F��H����W��^�W���u�u�d�`�j�}�G��H����W��^�D��e�d�e�d�g�l�[�ԜY����F�L�D��e�e�d�e�f�m�F��I����V��L����u�e�u�k�u�m�F��H����V��^�E��e�d�d�d�u�}�W���H���F�_�D��e�e�e�d�g�l�G��H����V�d��U��l�h�u�e�f�l�G��H����V��_�E��d�d�d�y�]�}�W��Y���V��_�E��d�e�d�d�f�m�F��I����FǻN��D���k�w�e�d�f�l�G��H����V��^�E��e�w�u�u�w�l�E��Y����W��^�E��d�d�e�e�g�m�G��H���F�_�H���e�d�d�e�g�l�G��I����V��^�D��y�_�u�u�f�}�I���I����W��_�D��e�e�d�d�g�m�G���Y���W��S�W��d�d�d�e�f�l�G��H����W��^�W���u�u�d�c�j�}�G��H����W��_�E��d�e�d�d�f�m�[�ԜY����F�L�D��e�e�d�e�f�l�F��I����V��L����u�d�u�k�u�m�F��H����V��_�D��e�d�d�e�u�}�W���H���F�_�D��e�d�e�e�f�l�F��I����V�d��U��e�h�u�e�f�l�G��H����V��_�D��d�d�d�y�]�}�W��Y���V��_�E��d�e�d�d�f�l�F��I����FǻN��G���k�w�e�d�f�l�G��H����W��_�D��d�w�u�u�w�l�D��Y����W��^�E��d�e�e�e�g�l�G��H���F�\�H���e�d�d�e�g�m�G��H����V��^�E��y�_�u�u�e�}�I���I����W��^�E��e�e�d�e�f�l�G���Y���W��S�W��d�d�d�d�g�l�F��H����W��_�W���u�u�d�b�j�}�G��H����V��_�D��e�d�e�e�g�l�[�ԜY����F�L�D��e�e�e�d�g�l�F��H����V��L����u�g�u�k�u�m�F��H����V��^�D��d�e�e�d�u�}�W���H���F�_�D��d�e�d�e�g�l�F��H����W�d��U��d�h�u�e�f�l�G��I����W��^�E��d�e�e�y�]�}�W��Y���V��_�E��d�d�e�e�g�m�F��H����FǻN��F���k�w�e�d�f�l�F��I����W��_�E��d�w�u�u�w�l�C��Y����W��^�D��e�d�e�d�g�l�G��I���F�]�H���e�d�d�e�g�m�G��H����W��_�E��y�_�u�u�d�}�I���I����W��_�E��e�d�e�e�g�l�F���Y���W��S�W��d�d�d�d�f�l�F��H����V��^�W���u�u�d�m�j�}�G��H����V��^�E��e�d�e�d�g�l�[�ԜY����
F�L�D��e�e�e�d�f�m�F��I����V��L����u�a�u�k�u�m�F��H����V��_�D��e�e�d�e�u�}�W���H���F�_�D��d�d�d�d�f�l�F��H����W�d��U��g�h�u�e�f�l�G��I����W��^�D��d�d�d�y�]�}�W��Y���V��_�E��e�e�d�e�g�l�F��I����FǻN��A���k�w�e�d�f�l�F��I����W��^�D��e�w�u�u�w�l�B��Y����W��^�E��d�e�e�d�f�l�G��I���F�Z�H���e�d�d�e�g�l�G��I����W��_�E��y�_�u�u�c�}�I���I����W��^�D��e�d�e�d�f�m�F���Y���W��S�W��d�d�d�d�g�m�G��H����W��^�W���u�u�d�l�j�}�G��H����W��^�D��e�d�d�d�g�l�[�ԜY����F�L�D��e�e�d�d�f�m�F��I����V��L����u�`�u�k�u�m�F��H����W��^�D��d�e�e�d�u�}�W���H���F�_�D��d�e�d�e�g�m�G��I����V�d��U��f�h�u�e�f�l�G��H����V��^�D��e�e�e�y�]�}�W��Y���V��_�E��e�e�d�e�g�l�G��I����FǻN��@���k�w�e�d�f�l�F��I����W��^�E��e�w�u�u�w�l�A��Y����W��^�D��e�d�e�d�f�l�G��H���F�[�H���e�d�d�e�g�l�G��I����W��^�D��y�_�u�u�b�}�I���I����W��_�E��e�d�e�d�f�m�F���Y���W��S�W��d�d�d�d�f�m�F��H����V��_�W���u�u�d�e�j�}�G��H����W��_�E��e�d�d�d�f�m�[�ԜY����F�L�D��e�e�d�d�g�l�F��I����V��L����u�c�u�k�u�m�F��H����W��_�D��e�d�d�d�u�}�W���H���F�_�D��d�d�d�d�f�l�F��I����W�d��U��a�h�u�e�f�l�G��I����W��_�E��e�d�e�y�]�}�W��Y���V��_�D��e�e�d�e�g�m�G��I����FǻN��C���k�w�e�d�f�l�G��I����V��_�D��d�w�u�u�w�l�@��Y����W��_�E��d�e�d�e�g�l�G��H���F�X�H���e�d�d�e�f�m�G��H����W��^�E��y�_�u�u�a�}�I���I����W��^�E��d�e�d�d�f�l�F���Y���W��S�W��d�d�d�e�g�l�F��I����W��^�W���u�u�d�d�j�}�G��H����V��_�E��d�e�d�d�f�m�[�ԜY����F�L�D��e�d�e�e�f�l�F��I����V��L����u�b�u�k�u�m�F��H����W��_�E��e�d�e�e�u�}�W���H���F�_�D��e�e�e�e�g�m�F��H����V�d��U��`�h�u�e�f�l�G��I����V��^�D��e�d�e�y�]�}�W��Y���V��_�D��d�d�e�d�g�m�G��H����FǻN��B���k�w�e�d�f�l�G��I����V��^�D��e�w�u�u�w�l�O��Y����W��_�E��d�e�d�e�f�m�F��I���F�Y�H���e�d�d�e�f�m�F��I����V��^�D��y�_�u�u�o�}�I���I����W��^�E��e�e�d�e�f�l�F���Y���W��S�W��d�d�d�e�g�l�G��I����W��_�W���u�u�d�g�j�}�G��H����V��_�D��e�d�e�d�g�l�[�ԜY���� F�L�D��e�d�e�d�f�l�G��I����V��L����u�m�u�k�u�m�F��H����V��_�E��d�d�e�e�u�}�W���H���F�_�D��e�d�e�d�g�m�F��H����W�d��U��c�h�u�e�f�l�G��I����W��^�D��d�e�e�y�]�}�W��Y���V��_�D��e�d�d�d�f�l�G��H����FǻN��M���k�w�e�d�f�l�G��I����V��^�D��d�w�u�u�w�l�N��Y����W��_�D��e�d�e�d�f�l�F��H���F�W�H���e�d�d�e�f�m�G��I����W��_�E��y�_�u�u�n�}�I���I����W��_�E��d�e�e�e�f�l�F���Y���W��S�W��d�d�d�e�f�l�G��I����V��_�W���u�u�d�f�j�}�G��H����V��_�D��e�d�e�e�g�m�[�ԜY����F�L�D��e�d�e�d�g�m�F��H����W��L����u�l�u�k�u�m�F��H����V��^�E��d�e�d�d�u�}�W���H���F�_�D��e�d�e�d�f�m�G��I����V�d��U��b�h�u�e�f�l�G��I����W��^�D��e�e�e�y�]�}�W��Y���V��_�D��d�d�e�e�f�m�G��I����FǻN��L���k�w�e�d�f�l�G��H����V��^�D��d�w�u�u�w�o�G��Y����W��_�D��e�d�e�d�g�l�F��H���F�^�H���e�d�d�e�f�m�F��H����V��_�E��y�_�u�u�g�}�I���I����W��_�D��d�d�e�d�f�m�F���Y���T��S�W��d�d�d�e�f�l�F��I����W��^�W���u�u�g�a�j�}�G��H����W��^�E��d�e�d�e�f�l�[�ԜY����F�L�D��e�d�d�e�g�l�G��H����V��L����u�e�u�k�u�m�F��H����V��^�D��d�d�e�e�u�}�W���K���F�_�D��e�e�e�e�f�m�G��I����W�d��U��m�h�u�e�f�l�G��H����V��^�E��e�d�e�y�]�}�W��Y���V��_�D��e�d�d�d�f�m�F��I����FǻN��D���k�w�e�d�f�l�G��H����V��_�D��e�w�u�u�w�o�F��Y����W��_�E��d�e�e�e�f�l�G��H���F�_�H���e�d�d�e�f�l�G��I����W��_�E��y�_�u�u�f�}�I���I����W��^�D��e�d�d�d�g�m�G���Y���T��S�W��d�d�d�e�g�l�F��I����W��^�W���u�u�g�`�j�}�G��H����W��^�E��e�d�d�d�g�m�[�ԜY����F�L�D��e�d�d�d�g�m�F��H����W��L����u�d�u�k�u�m�F��H����V��^�D��e�e�d�e�u�}�W���K���F�_�D��e�e�e�d�g�m�F��H����V�d��U��l�h�u�e�f�l�G��H����W��_�E��d�e�d�y�]�}�W��Y���V��_�D��d�e�d�e�g�m�G��H����FǻN��G���k�w�e�d�f�l�G��H����W��_�E��d�w�u�u�w�o�E��Y����W��_�E��e�e�e�d�f�l�F��H���F�\�H���e�d�d�e�f�l�F��H����W��_�D��y�_�u�u�e�}�I���I����W��^�D��d�e�d�d�g�m�G���Y���T��S�W��d�d�d�e�f�m�G��H����W��^�W���u�u�g�c�j�}�G��H����W��^�D��d�d�e�e�g�l�[�ԜY����F�L�D��e�d�d�e�f�m�G��H����W��L����u�g�u�k�u�m�F��H����V��_�E��d�d�d�d�u�}�W���K���F�_�D��e�d�e�d�g�m�G��I����W�d��U��e�h�u�e�f�l�G��H����V��_�E��e�d�e�y�]�}�W��Y���V��_�D��e�e�e�d�g�m�F��I����FǻN��F���k�w�e�d�f�l�G��H����W��^�E��d�w�u�u�w�o�D��Y����W��_�D��e�d�e�e�f�m�F��H���F�]�H���e�d�d�e�f�l�G��H����V��^�D��y�_�u�u�d�}�I���I����W��_�E��e�e�e�d�g�l�F���Y���T��S�W��d�d�d�e�f�m�F��H����W��_�W���u�u�g�b�j�}�G��H����W��^�D��e�e�e�d�g�l�[�ԜY����F�L�D��e�d�d�d�f�l�F��H����V��L����u�f�u�k�u�m�F��H����V��_�E��d�e�d�e�u�}�W���K���F�_�D��e�d�d�e�g�l�G��H����W�d��U��d�h�u�e�f�l�G��H����V��^�E��d�e�e�y�]�}�W��Y���V��_�D��d�e�d�e�f�l�G��H����FǻN��A���k�w�e�d�f�l�G��H����W��_�E��e�w�u�u�w�o�C��Y����W��_�D��d�d�d�e�f�m�G��H���F�Z�H���e�d�d�e�f�m�G��I����W��_�E��y�_�u�u�c�}�I���I����W��^�E��d�d�d�d�f�m�F���Y���T��S�W��d�d�d�d�g�m�F��H����V��^�W���u�u�g�m�j�}�G��H����V��_�D��d�e�e�d�g�l�[�ԜY����
F�L�D��e�d�e�e�f�m�G��I����W��L����u�`�u�k�u�m�F��H����W��^�D��d�e�e�d�u�}�W���K���F�_�D��d�e�d�e�f�l�F��I����V�d��U��g�h�u�e�f�l�G��I����W��_�E��e�d�e�y�]�}�W��Y���V��_�D��e�d�e�d�g�m�F��I����FǻN��@���k�w�e�d�f�l�F��H����V��_�E��d�w�u�u�w�o�B��Y����W��_�E��d�d�d�d�f�m�F��H���F�[�H���e�d�d�e�f�m�F��H����V��_�D��y�_�u�u�b�}�I���I����W��^�E��e�e�e�e�g�l�G���Y���T��S�W��d�d�d�d�g�m�G��I����W��^�W���u�u�g�l�j�}�G��H����V��_�E��d�d�d�d�f�l�[�ԜY����F�L�D��e�d�e�d�f�l�G��I����V��L����u�c�u�k�u�m�F��H����W��^�E��d�e�e�d�u�}�W���K���F�_�D��d�e�d�d�f�m�F��I����W�d��U��f�h�u�e�f�l�G��I����V��^�D��e�d�e�y�]�}�W��Y���V��_�D��d�d�d�d�f�m�F��I����FǻN��C���k�w�e�d�f�l�F��H����V��_�D��d�w�u�u�w�o�A��Y����W��_�D��e�e�e�d�f�l�G��I���F�X�H���e�d�d�e�f�m�G��I����V��^�D��y�_�u�u�a�}�I���I����W��_�D��e�d�e�d�g�l�G���Y���T��S�W��d�d�d�d�f�m�G��I����W��^�W���u�u�g�e�j�}�G��H����V��_�E��d�d�d�e�f�l�[�ԜY����F�L�D��e�d�e�e�g�m�F��I����V��L����u�b�u�k�u�m�F��H����W��^�D��d�d�d�e�u�}�W���K���F�_�D��d�d�d�e�g�m�F��I����V�d��U��a�h�u�e�f�l�G��I����W��_�D��e�d�d�y�]�}�W��Y���V��_�D��e�d�d�e�g�m�F��H����FǻN��B���k�w�e�d�f�l�F��I����W��_�E��e�w�u�u�w�o�@��Y����W��_�D��d�e�e�d�f�l�F��I���F�Y�H���e�d�d�e�f�m�F��H����V��_�D��y�_�u�u�`�}�I���I����W��_�D��d�e�e�e�g�l�F���Y���T��S�W��d�d�d�d�f�m�F��H����V��_�W���u�u�g�d�j�}�G��H����V��^�D��d�d�e�d�f�m�[�ԜY����F�L�D��e�d�e�d�g�m�G��I����V��L����u�m�u�k�u�m�F��H����W��_�E��d�d�e�e�u�}�W���K���F�_�D��d�d�d�e�g�l�F��H����V�d��U��`�h�u�e�f�l�G��I����V��^�E��e�e�e�y�]�}�W��Y���V��_�D��e�e�e�d�f�m�G��H����FǻN��M���k�w�e�d�f�l�F��I����W��^�E��d�w�u�u�w�o�O��Y����W��_�E��d�e�d�d�g�m�G��I���F�V�H���e�d�d�e�f�l�G��H����V��^�E��y�_�u�u�n�}�I���I����W��^�D��e�d�d�d�g�m�F���Y���T��S�W��d�d�d�d�g�l�G��H����V��_�W���u�u�g�g�j�}�G��H����W��^�D��e�d�d�d�f�m�[�ԜY���� F�L�D��e�d�d�e�g�l�F��H����V��L����u�l�u�k�u�m�F��H����W��_�D��e�e�d�e�u�}�W���K���F�_�D��d�e�d�d�g�l�G��H����V�d��U��c�h�u�e�f�l�G��H����W��_�E��d�e�e�y�]�}�W��Y���V��_�D��d�e�d�e�g�l�G��H����FǻN��L���k�w�e�d�f�l�F��I����V��^�E��d�w�u�u�w�o�N��Y����W��_�E��e�d�d�e�f�l�F��I���F�^�H���e�d�d�e�f�l�F��I����V��^�E��y�_�u�u�g�}�I���I����W��^�D��d�e�e�e�g�m�G���Y���U��S�W��d�d�d�d�g�l�G��I����V��_�W���u�u�f�f�j�}�G��H����W��^�D��e�e�d�e�g�l�[�ԜY����F�L�D��e�d�d�d�f�m�F��I����V��L����u�e�u�k�u�m�F��H����W��^�E��e�d�d�e�u�}�W���J���F�_�D��d�e�d�d�f�m�F��H����W�d��U��b�h�u�e�f�l�G��H����W��_�D��e�e�d�y�]�}�W��Y���V��_�D��e�e�e�e�g�l�G��H����FǻN��E���k�w�e�d�f�l�F��I����W��^�E��d�w�u�u�w�n�G��Y����W��_�D��e�d�e�d�g�l�F��I���F�_�H���e�d�d�e�f�l�G��H����W��^�D��y�_�u�u�f�}�I���I����W��_�E��d�e�e�d�g�m�G���Y���U��S�W��d�d�d�d�f�l�F��H����W��_�W���u�u�f�a�j�}�G��H����W��_�E��d�e�d�d�g�l�[�ԜY����F�L�D��e�d�d�e�f�l�G��I����V��L����u�d�u�k�u�m�F��H����W��^�E��e�d�d�e�u�}�W���J���F�_�D��d�d�e�e�f�l�G��H����V�d��U��m�h�u�e�f�l�G��H����V��^�D��d�d�e�y�]�}�W��Y���V��_�D��d�e�d�d�f�l�F��I����FǻN��G���k�w�e�d�f�l�F��I����W��^�D��d�w�u�u�w�n�F��Y����W��_�D��d�d�d�e�f�l�F��I���F�\�H���e�d�d�e�f�l�F��I����V��^�D��y�_�u�u�e�}�I���I����W��_�E��e�d�e�e�g�l�F���Y���U��S�W��d�d�d�d�f�l�F��H����V��^�W���u�u�f�`�j�}�G��H����W��_�E��e�e�e�d�f�m�[�ԜY����F�L�D��e�d�d�d�f�m�G��H����V��L����u�g�u�k�u�m�F��I����V��^�E��d�e�d�e�u�}�W���J���F�_�D��e�e�e�e�f�l�F��H����W�d��U��l�h�u�e�f�l�F��I����W��_�D��e�e�d�y�]�}�W��Y���V��_�E��e�e�e�d�f�l�F��H����FǻN��F���k�w�e�d�f�m�G��I����V��^�D��d�w�u�u�w�n�E��Y����W��^�E��e�e�e�d�g�m�G��I���F�]�H���e�d�d�d�g�m�G��I����V��_�D��y�_�u�u�d�}�I���I����V��^�D��e�d�e�d�g�l�F���Y���U��S�W��d�d�e�e�g�m�F��H����W��_�W���u�u�f�c�j�}�G��H����V��_�E��d�d�e�e�g�m�[�ԜY����F�L�D��d�e�e�e�f�l�F��I����V��L����u�f�u�k�u�m�F��I����W��_�D��e�d�e�e�u�}�W���J���F�_�D��e�e�d�e�f�m�G��I����V�d��U��e�h�u�e�f�l�F��I����V��^�D��e�e�e�y�]�}�W��Y���V��_�E��e�e�d�e�g�l�G��H����FǻN��A���k�w�e�d�f�m�G��H����V��_�E��d�w�u�u�w�n�D��Y����W��^�E��e�d�e�d�g�l�G��H���F�Z�H���e�d�d�d�g�m�G��H����W��_�D��y�_�u�u�c�}�I���I����V��^�D��e�e�d�e�g�m�F���Y���U��S�W��d�d�e�e�g�l�F��H����V��_�W���u�u�f�b�j�}�G��H����V��_�D��d�d�d�e�g�l�[�ԜY����F�L�D��d�e�e�d�g�m�G��I����V��L����u�a�u�k�u�m�F��I����V��^�E��d�d�e�d�u�}�W���J���F�_�D��e�e�e�d�g�m�G��H����V�d��U��d�h�u�e�f�l�F��I����V��_�D��e�e�e�y�]�}�W��Y���V��_�E��d�e�d�e�f�l�F��I����FǻN��@���k�w�e�d�f�m�G��I����W��_�D��e�w�u�u�w�n�C��Y����W��^�E��e�e�d�d�g�m�F��H���F�[�H���e�d�d�d�g�m�F��H����W��^�E��y�_�u�u�b�}�I���I����V��^�D��e�d�e�d�f�m�F���Y���U��S�W��d�d�e�e�g�m�F��I����V��^�W���u�u�f�m�j�}�G��H����V��^�E��d�d�e�e�g�l�[�ԜY����
F�L�D��d�e�e�d�g�l�G��I����V��L����u�c�u�k�u�m�F��I����W��_�D��e�e�d�d�u�}�W���J���F�_�D��e�e�d�d�f�m�F��H����V�d��U��g�h�u�e�f�l�F��I����W��^�D��e�d�d�y�]�}�W��Y���V��_�E��d�d�e�e�g�l�F��H����FǻN��C���k�w�e�d�f�m�G��H����W��^�E��d�w�u�u�w�n�B��Y����W��^�E��e�d�d�d�g�m�F��I���F�X�H���e�d�d�d�g�m�F��I����V��_�D��y�_�u�u�a�}�I���I����V��^�D��d�e�e�e�f�l�F���Y���U��S�W��d�d�e�e�f�m�G��I����V��_�W���u�u�f�l�j�}�G��H����V��^�D��d�e�e�d�f�m�[�ԜY����F�L�D��d�e�e�e�g�l�G��H����V��L����u�b�u�k�u�m�F��I����V��^�E��e�e�d�e�u�}�W���J���F�_�D��e�d�e�d�g�l�F��H����V�d��U��f�h�u�e�f�l�F��I����W��_�E��e�d�e�y�]�}�W��Y���V��_�E��e�d�e�e�f�m�F��H����FǻN��B���k�w�e�d�f�m�G��I����V��_�E��e�w�u�u�w�n�A��Y����W��^�D��d�e�e�d�g�l�G��I���F�Y�H���e�d�d�d�g�m�G��H����V��^�D��y�_�u�u�`�}�I���I����V��_�D��d�d�d�d�g�m�G���Y���U��S�W��d�d�e�e�f�l�G��I����V��^�W���u�u�f�e�j�}�G��H����V��^�E��e�e�e�d�g�m�[�ԜY����F�L�D��d�e�e�e�g�m�G��H����W��L����u�m�u�k�u�m�F��I����W��_�D��d�e�d�d�u�}�W���J���F�_�D��e�d�d�d�f�l�F��I����W�d��U��a�h�u�e�f�l�F��I����V��^�E��e�e�d�y�]�}�W��Y���V��_�E��e�d�d�d�g�l�F��I����FǻN��M���k�w�e�d�f�m�G��H����V��_�D��d�w�u�u�w�n�@��Y����W��^�D��d�d�e�e�g�l�F��H���F�V�H���e�d�d�d�g�m�G��H����W��_�D��y�_�u�u�o�}�I���I����V��_�E��d�e�e�d�f�l�G���Y���U��S�W��d�d�e�e�f�m�G��H����V��^�W���u�u�f�d�j�}�G��H����V��^�D��e�e�d�d�g�l�[�ԜY����F�L�D��d�e�e�d�g�m�G��H����V��L����u�l�u�k�u�m�F��I����V��^�D��e�e�e�e�u�}�W���J���F�_�D��e�d�e�e�g�m�G��I����V�d��U��`�h�u�e�f�l�F��I����W��^�E��e�e�e�y�]�}�W��Y���V��_�E��d�d�d�d�f�m�G��H����FǻN��L���k�w�e�d�f�m�G��I����V��^�E��d�w�u�u�w�n�O��Y����W��^�D��d�e�d�e�g�m�G��H���F�W�H���e�d�d�d�g�m�F��I����W��^�E��y�_�u�u�g�}�I���I����V��_�E��d�e�d�d�g�l�F���Y���R��S�W��d�d�e�e�f�l�G��H����V��_�W���u�u�a�g�j�}�G��H����V��^�E��d�d�e�e�f�m�[�ԜY���� F�L�D��d�e�e�d�g�l�F��I����V��L����u�e�u�k�u�m�F��I����W��^�E��e�d�d�e�u�}�W���M���F�_�D��e�d�d�e�f�m�F��I����W�d��U��c�h�u�e�f�l�F��I����W��_�E��d�d�d�y�]�}�W��Y���V��_�E��d�d�e�d�f�l�G��H����FǻN��E���k�w�e�d�f�m�G��H����W��_�D��d�w�u�u�w�i�N��Y����W��^�D��d�d�d�d�g�l�G��I���F�_�H���e�d�d�d�g�l�G��I����V��^�E��y�_�u�u�f�}�I���I����V��^�E��d�d�d�e�g�l�G���Y���R��S�W��d�d�e�e�g�m�F��H����V��_�W���u�u�a�f�j�}�G��H����W��^�E��e�d�d�e�g�l�[�ԜY����F�L�D��d�e�d�e�g�l�F��I����V��L����u�d�u�k�u�m�F��I����V��_�D��e�d�e�e�u�}�W���M���F�_�D��e�e�e�e�g�m�G��I����V�d��U��b�h�u�e�f�l�F��H����V��_�E��d�d�e�y�]�}�W��Y���V��_�E��e�d�e�d�g�l�G��I����FǻN��D���k�w�e�d�f�m�G��I����W��_�D��d�w�u�u�w�i�G��Y����W��^�E��e�e�d�e�g�m�G��H���F�\�H���e�d�d�d�g�l�G��H����W��_�D��y�_�u�u�e�}�I���I����V��^�E��d�d�d�e�f�m�G���Y���R��S�W��d�d�e�e�g�l�F��I����W��_�W���u�u�a�a�j�}�G��H����W��^�D��d�d�e�e�f�m�[�ԜY����F�L�D��d�e�d�e�f�m�F��I����V��L����u�g�u�k�u�m�F��I����W��^�D��d�d�e�d�u�}�W���M���F�_�D��e�e�d�e�f�m�F��I����V�d��U��m�h�u�e�f�l�F��H����V��^�E��d�e�d�y�]�}�W��Y���V��_�E��e�d�d�d�g�m�G��H����FǻN��F���k�w�e�d�f�m�G��I����W��^�D��d�w�u�u�w�i�F��Y����W��^�E��e�d�d�e�f�l�F��I���F�]�H���e�d�d�d�g�l�F��H����W��_�D��y�_�u�u�d�}�I���I����V��^�E��e�e�d�e�f�m�F���Y���R��S�W��d�d�e�e�g�m�F��I����W��^�W���u�u�a�`�j�}�G��H����W��_�E��e�e�d�e�g�l�[�ԜY����F�L�D��d�e�d�d�f�m�F��H����W��L����u�f�u�k�u�m�F��I����V��_�D��d�d�d�d�u�}�W���M���F�_�D��e�e�e�d�g�l�G��H����V�d��U��l�h�u�e�f�l�F��H����W��^�E��e�e�d�y�]�}�W��Y���V��_�E��d�d�d�d�f�m�G��I����FǻN��A���k�w�e�d�f�m�G��H����W��_�E��d�w�u�u�w�i�E��Y����W��^�E��e�e�d�d�g�m�F��I���F�Z�H���e�d�d�d�g�l�F��I����V��^�D��y�_�u�u�c�}�I���I����V��^�E��e�e�e�e�f�m�G���Y���R��S�W��d�d�e�e�g�l�F��I����W��^�W���u�u�a�c�j�}�G��H����W��_�D��e�e�e�e�f�l�[�ԜY����F�L�D��d�e�d�d�f�l�F��I����V��L����u�a�u�k�u�m�F��I����W��^�E��d�d�e�d�u�}�W���M���F�_�D��e�e�d�d�f�l�G��I����V�d��U��e�h�u�e�f�l�F��H����W��^�E��d�e�d�y�]�}�W��Y���V��_�E��e�e�e�d�f�m�F��I����FǻN��@���k�w�e�d�f�m�G��I����W��^�E��e�w�u�u�w�i�D��Y����W��^�D��e�d�d�d�f�l�G��I���F�[�H���e�d�d�d�g�l�G��I����W��^�E��y�_�u�u�b�}�I���I����V��_�E��e�e�e�d�g�m�G���Y���R��S�W��d�d�e�e�f�m�G��I����W��_�W���u�u�a�b�j�}�G��H����W��_�E��e�d�d�d�g�l�[�ԜY����F�L�D��d�e�d�e�f�l�F��H����W��L����u�`�u�k�u�m�F��I����V��_�E��d�e�d�d�u�}�W���M���F�_�D��e�d�e�d�g�l�F��H����V�d��U��d�h�u�e�f�l�F��H����V��^�D��d�d�e�y�]�}�W��Y���V��_�E��e�e�e�d�f�l�F��I����FǻN��C���k�w�e�d�f�m�G��H����W��_�D��d�w�u�u�w�i�C��Y����W��^�D��d�d�e�e�g�m�F��I���F�X�H���e�d�d�d�g�l�G��H����W��^�E��y�_�u�u�a�}�I���I����V��_�D��e�e�d�e�f�l�G���Y���R��S�W��d�d�e�e�f�l�G��I����W��_�W���u�u�a�m�j�}�G��H����W��_�D��d�e�d�d�g�m�[�ԜY����
F�L�D��d�e�d�e�f�m�F��H����W��L����u�b�u�k�u�m�F��I����W��^�E��e�d�e�d�u�}�W���M���F�_�D��e�d�d�d�f�l�F��I����V�d��U��g�h�u�e�f�l�F��H����V��^�D��e�d�e�y�]�}�W��Y���V��_�E��d�e�d�d�f�l�F��H����FǻN��B���k�w�e�d�f�m�G��I����W��_�D��e�w�u�u�w�i�B��Y����W��^�D��d�e�e�e�g�m�G��H���F�Y�H���e�d�d�d�g�l�F��H����W��_�D��y�_�u�u�`�}�I���I����V��_�D��e�e�d�e�g�m�F���Y���R��S�W��d�d�e�e�f�m�G��I����V��^�W���u�u�a�l�j�}�G��H����W��_�E��e�d�d�d�g�l�[�ԜY����F�L�D��d�e�d�d�f�m�F��H����W��L����u�m�u�k�u�m�F��I����V��_�E��d�d�e�d�u�}�W���M���F�_�D��e�d�d�e�g�l�F��H����V�d��U��f�h�u�e�f�l�F��H����W��^�D��e�d�e�y�]�}�W��Y���V��_�E��d�e�d�d�f�l�G��I����FǻN��M���k�w�e�d�f�m�G��H����W��^�D��d�w�u�u�w�i�A��Y����W��^�D��d�e�d�d�f�m�G��H���F�V�H���e�d�d�d�g�l�F��I����W��_�D��y�_�u�u�o�}�I���I����V��_�D��e�e�e�e�f�l�F���Y���R��S�W��d�d�e�e�f�l�G��I����V��_�W���u�u�a�e�j�}�G��H����W��_�D��e�e�d�e�f�l�[�ԜY����F�L�D��d�e�d�d�f�l�F��I����W��L����u�l�u�k�u�m�F��I����V��^�E��e�e�d�e�u�}�W���M���F�_�D��d�e�e�e�f�l�G��I����V�d��U��a�h�u�e�f�l�F��I����W��^�D��e�d�e�y�]�}�W��Y���V��_�E��e�e�e�d�f�m�G��H����FǻN��L���k�w�e�d�f�m�F��I����W��_�D��d�w�u�u�w�i�@��Y����W��^�E��d�d�d�d�f�l�G��I���F�W�H���e�d�d�d�g�m�G��I����V��_�E��y�_�u�u�n�}�I���I����V��^�D��e�e�d�e�g�m�F���Y���S��S�W��d�d�e�d�g�m�F��I����V��_�W���u�u�`�d�j�}�G��H����V��_�E��e�e�e�d�f�l�[�ԜY����F�L�D��d�e�e�e�f�l�F��H����V��L����u�e�u�k�u�m�F��I����W��_�D��e�e�e�e�u�}�W���L���F�_�D��d�e�d�e�g�l�G��I����W�d��U���`�h�u�e�f�l�F��I����V��^�D��e�e�d�y�]�}�W��Y���V��_�E��e�e�e�d�g�l�G��I����FǻN��E���k�w�e�d�f�m�F��H����W��^�D��d�w�u�u�w�h�O��Y����W��^�E��e�e�d�e�f�l�G��H���F�^�H���e�d�d�d�g�m�G��H����V��_�D��y�_�u�u�f�}�I���I����V��^�D��e�e�e�d�g�l�F���Y���S��S�W��d�d�e�d�g�l�F��I����V��^�W���u�u�`�g�j�}�G��H����V��_�D��d�d�d�e�g�m�[�ԜY���� F�L�D��d�e�e�d�g�m�F��I����W��L����u�d�u�k�u�m�F��I����V��^�D��d�d�e�e�u�}�W���L���F�_�D��d�e�e�e�f�m�F��I����W�d��U���c�h�u�e�f�l�F��I����V��^�E��d�e�e�y�]�}�W��Y���V��_�E��d�e�d�d�g�l�F��H����FǻN��D���k�w�e�d�f�m�F��I����W��_�D��e�w�u�u�w�h�N��Y����W��^�E��e�d�d�d�f�l�G��I���F�\�H���e�d�d�d�g�m�F��H����W��^�D��y�_�u�u�e�}�I���I����V��^�D��d�d�e�d�g�l�G���Y���S��S�W��d�d�e�d�g�m�F��H����W��_�W���u�u�`�f�j�}�G��H����V��^�E��e�d�d�e�f�m�[�ԜY����F�L�D��d�e�e�d�g�m�F��I����V��L����u�g�u�k�u�m�F��I����W��_�E��d�d�d�e�u�}�W���L���F�_�D��d�e�d�d�g�m�G��H����W�d��U���b�h�u�e�f�l�F��I����W��_�D��e�d�e�y�]�}�W��Y���V��_�E��d�e�d�d�f�l�G��I����FǻN��G���k�w�e�d�f�m�F��H����W��^�E��e�w�u�u�w�h�G��Y����W��^�E��e�e�d�e�f�l�F��I���F�]�H���e�d�d�d�g�m�F��I����V��^�D��y�_�u�u�d�}�I���I����V��^�D��d�d�e�e�f�l�G���Y���S��S�W��d�d�e�d�g�l�F��H����V��^�W���u�u�`�a�j�}�G��H����V��^�E��d�d�e�d�g�l�[�ԜY����F�L�D��d�e�e�e�g�l�G��H����V��L����u�f�u�k�u�m�F��I����V��^�E��d�d�e�e�u�}�W���L���F�_�D��d�d�e�d�f�m�F��H����V�d��U���m�h�u�e�f�l�F��I����W��^�E��e�e�d�y�]�}�W��Y���V��_�E��e�d�e�d�f�m�G��I����FǻN��A���k�w�e�d�f�m�F��I����V��_�E��e�w�u�u�w�h�F��Y����W��^�D��e�d�e�d�f�l�G��I���F�Z�H���e�d�d�d�g�m�G��I����V��^�E��y�_�u�u�c�}�I���I����V��_�D��d�e�d�d�f�m�F���Y���S��S�W��d�d�e�d�f�l�G��H����V��^�W���u�u�`�`�j�}�G��H����V��^�D��d�d�d�d�g�m�[�ԜY����F�L�D��d�e�e�e�g�l�G��I����V��L����u�a�u�k�u�m�F��I����W��^�D��e�e�e�d�u�}�W���L���F�_�D��d�d�d�d�g�l�F��H����V�d��U���l�h�u�e�f�l�F��I����V��^�E��e�e�d�y�]�}�W��Y���V��_�E��e�d�e�d�g�l�F��H����FǻN��@���k�w�e�d�f�m�F��H����V��_�E��e�w�u�u�w�h�E��Y����W��^�D��d�e�e�d�f�m�G��H���F�[�H���e�d�d�d�g�m�G��H����V��^�D��y�_�u�u�b�}�I���I����V��_�D��d�d�e�e�g�l�G���Y���S��S�W��d�d�e�d�f�m�G��I����W��^�W���u�u�`�c�j�}�G��H����V��^�E��e�e�e�e�f�m�[�ԜY����F�L�D��d�e�e�d�g�m�G��H����V��L����u�`�u�k�u�m�F��I����V��_�E��e�d�e�d�u�}�W���L���F�_�D��d�d�e�d�f�l�F��H����V�d��U���e�h�u�e�f�l�F��I����V��_�D��d�d�d�y�]�}�W��Y���V��_�E��d�d�d�e�f�l�F��H����FǻN��C���k�w�e�d�f�m�F��I����W��^�E��e�w�u�u�w�h�D��Y����W��^�D��d�d�e�e�g�m�F��I���F�X�H���e�d�d�d�g�m�F��H����W��_�E��y�_�u�u�a�}�I���I����V��_�E��d�e�e�d�g�l�G���Y���S��S�W��d�d�e�d�f�l�G��I����W��_�W���u�u�`�b�j�}�G��H����V��^�D��e�e�d�d�g�l�[�ԜY����F�L�D��d�e�e�d�g�m�G��H����W��L����u�c�u�k�u�m�F��I����W��^�D��e�e�e�e�u�}�W���L���F�_�D��d�d�d�e�g�m�F��H����W�d��U���d�h�u�e�f�l�F��I����V��^�D��e�d�d�y�]�}�W��Y���V��_�E��d�d�d�e�g�l�F��H����FǻN��B���k�w�e�d�f�m�F��H����W��_�E��d�w�u�u�w�h�C��Y����W��^�D��d�e�d�d�f�l�G��I���F�Y�H���e�d�d�d�g�m�F��H����V��_�D��y�_�u�u�`�}�I���I����V��^�E��e�d�e�e�g�m�F���Y���S��S�W��d�d�e�d�g�m�G��H����V��^�W���u�u�`�m�j�}�G��H����W��^�E��e�e�e�d�f�m�[�ԜY����
F�L�D��d�e�d�e�g�l�G��H����W��L����u�m�u�k�u�m�F��I����V��_�E��e�e�d�e�u�}�W���L���F�_�D��d�e�e�e�f�m�F��H����W�d��U���g�h�u�e�f�l�F��H����W��_�E��d�d�e�y�]�}�W��Y���V��_�E��e�d�e�e�f�l�G��H����FǻN��M���k�w�e�d�f�m�F��I����V��^�E��d�w�u�u�w�h�B��Y����W��^�E��d�d�e�d�g�m�G��H���F�V�H���e�d�d�d�g�l�G��I����V��^�E��y�_�u�u�o�}�I���I����V��^�E��e�e�d�d�g�l�G���Y���S��S�W��d�d�e�d�g�l�G��H����V��_�W���u�u�`�l�j�}�G��H����W��^�D��d�e�e�e�g�l�[�ԜY����F�L�D��d�e�d�e�g�l�F��I����W��L����u�l�u�k�u�m�F��I����W��^�D��e�d�e�e�u�}�W���L���F�_�D��d�e�d�e�f�l�F��H����V�d��U���f�h�u�e�f�l�F��H����W��_�E��d�e�e�y�]�}�W��Y���V��_�E��e�d�e�e�g�m�G��H����FǻN��L���k�w�e�d�f�m�F��H����V��^�D��d�w�u�u�w�h�A��Y����W��^�E��e�e�e�d�g�m�G��I���F�W�H���e�d�d�d�g�l�F��I����W��^�E��y�_�u�u�n�}�I���I����V��^�E��e�e�d�d�f�m�F���Y���S��S�W��d�d�e�d�g�m�F��I����W��^�W���u�u�c�e�j�}�G��H����W��^�E��e�d�e�d�g�m�[�ԜY����F�L�D��d�e�d�d�g�l�F��I����W��L����u�e�u�k�u�m�F��I����V��_�D��e�d�d�e�u�}�W���O���F�_�D��d�e�e�e�g�l�G��H����W�d��U��a�h�u�e�f�l�F��H����V��^�D��e�d�d�y�]�}�W��Y���V��_�E��d�d�e�d�g�m�G��I����FǻN��E���k�w�e�d�f�m�F��I����W��^�E��e�w�u�u�w�k�@��Y����W��^�E��e�e�d�e�g�m�G��H���F�^�H���e�d�d�d�g�l�F��H����W��_�D��y�_�u�u�g�}�I���I����V��^�E��d�d�e�e�g�l�F���Y���P��S�W��d�d�e�d�g�l�F��H����V��^�W���u�u�c�d�j�}�G��H����W��^�E��d�d�d�e�g�l�[�ԜY����F�L�D��d�e�d�d�f�m�F��I����W��L����u�d�u�k�u�m�F��I����W��^�E��e�d�e�e�u�}�W���O���F�_�D��d�e�d�e�f�m�F��I����W�d��U��`�h�u�e�f�l�F��H����V��^�E��d�d�e�y�]�}�W��Y���V��_�E��d�d�d�d�f�m�F��I����FǻN��D���k�w�e�d�f�m�F��I����V��^�D��d�w�u�u�w�k�O��Y����W��^�D��e�d�e�d�g�m�G��I���F�_�H���e�d�d�d�g�l�G��H����V��^�D��y�_�u�u�e�}�I���I����V��_�E��d�d�d�d�g�m�G���Y���P��S�W��d�d�e�d�f�m�F��H����W��_�W���u�u�c�g�j�}�G��H����W��^�D��e�e�d�d�f�l�[�ԜY���� F�L�D��d�e�d�e�f�m�G��I����V��L����u�g�u�k�u�m�F��I����V��^�E��e�e�e�e�u�}�W���O���F�_�D��d�d�e�d�g�l�F��H����V�d��U��c�h�u�e�f�l�F��H����V��_�D��e�e�d�y�]�}�W��Y���V��_�E��e�d�d�e�f�l�G��I����FǻN��G���k�w�e�d�f�m�F��H����W��^�D��e�w�u�u�w�k�N��Y����W��^�D��e�e�d�d�g�m�G��I���F�]�H���e�d�d�d�g�l�G��I����V��_�D��y�_�u�u�d�}�I���I����V��_�E��d�e�e�d�g�m�G���Y���P��S�W��d�d�e�d�f�l�F��I����W��^�W���u�u�c�f�j�}�G��H����W��_�E��d�e�d�d�g�l�[�ԜY����F�L�D��d�e�d�e�f�l�G��H����V��L����u�f�u�k�u�m�F��I����W��_�D��e�e�e�d�u�}�W���O���F�_�D��d�d�d�d�f�m�G��I����V�d��U��b�h�u�e�f�l�F��H����W��_�D��d�e�d�y�]�}�W��Y���V��_�E��d�e�e�e�f�m�F��H����FǻN��F���k�w�e�d�f�m�F��I����V��^�E��d�w�u�u�w�k�G��Y����W��^�D��e�d�e�d�f�l�G��I���F�Z�H���e�d�d�d�g�l�F��I����V��^�D��y�_�u�u�c�}�I���I����V��_�E��e�e�d�d�g�m�G���Y���P��S�W��d�d�e�d�f�m�F��H����W��_�W���u�u�c�a�j�}�G��H����W��_�D��d�d�d�e�g�l�[�ԜY����F�L�D��d�e�d�d�f�l�F��H����V��L����u�a�u�k�u�m�F��I����V��^�D��d�d�d�e�u�}�W���O���F�_�D��d�d�e�d�f�l�G��I����W�d��U��m�h�u�e�f�l�F��H����W��_�D��e�d�e�y�]�}�W��Y���V��_�E��d�e�e�d�f�m�G��I����FǻN��@���k�w�e�d�f�m�F��H����W��^�E��d�w�u�u�w�k�F��Y����W��^�D��e�d�d�d�f�l�G��H���F�[�H���e�d�d�d�g�l�F��I����V��^�D��y�_�u�u�b�}�I���I����V��_�E��e�e�d�d�f�l�G���Y���P��S�W��d�d�e�d�f�l�G��I����V��^�W���u�u�c�`�j�}�G��H����W��_�E��d�d�e�e�g�m�[�ԜY����F�L�D��d�e�d�d�f�l�F��H����V��L����u�`�u�k�u�m�F��I����W��_�D��e�d�d�e�u�}�W���O���F�_�D��d�d�d�d�g�m�G��I����V�d��U��l�h�u�e�f�l�F��I����V��^�D��d�e�e�y�]�}�W��Y���V��_�D��e�e�e�d�g�l�G��I����FǻN��C���k�w�e�d�f�m�G��I����V��^�E��e�w�u�u�w�k�E��Y����W��_�E��e�e�d�d�f�l�F��I���F�X�H���e�d�d�d�f�m�G��H����V��^�E��y�_�u�u�a�}�I���I����V��^�E��d�d�e�d�g�m�G���Y���P��S�W��d�d�e�e�g�m�F��I����W��_�W���u�u�c�c�j�}�G��H����V��^�D��e�e�e�e�g�m�[�ԜY����F�L�D��d�d�e�e�g�l�G��H����W��L����u�c�u�k�u�m�F��I����V��^�D��e�e�d�d�u�}�W���O���F�_�D��e�e�e�d�f�m�G��H����V�d��U��e�h�u�e�f�l�F��I����V��_�E��e�e�e�y�]�}�W��Y���V��_�D��e�d�e�e�f�m�G��I����FǻN��B���k�w�e�d�f�m�G��I����W��_�E��e�w�u�u�w�k�D��Y����W��_�E��e�e�e�d�g�l�F��H���F�Y�H���e�d�d�d�f�m�G��H����W��_�D��y�_�u�u�`�}�I���I����V��^�D��e�d�d�d�g�l�G���Y���P��S�W��d�d�e�e�g�m�F��I����V��^�W���u�u�c�b�j�}�G��H����V��_�D��e�e�e�d�g�m�[�ԜY����F�L�D��d�d�e�e�f�l�F��I����W��L����u�b�u�k�u�m�F��I����V��_�E��d�e�d�d�u�}�W���O���F�_�D��e�e�d�e�g�m�G��H����V�d��U��d�h�u�e�f�l�F��I����V��^�D��e�e�e�y�]�}�W��Y���V��_�D��e�e�e�d�g�l�F��H����FǻN��M���k�w�e�d�f�m�G��H����W��^�E��e�w�u�u�w�k�C��Y����W��_�E��e�d�e�d�g�m�G��I���F�V�H���e�d�d�d�f�m�G��H����V��_�D��y�_�u�u�o�}�I���I����V��^�E��d�e�e�d�f�l�F���Y���P��S�W��d�d�e�e�g�l�F��H����W��_�W���u�u�c�m�j�}�G��H����V��^�E��d�e�d�e�f�m�[�ԜY����
F�L�D��d�d�e�e�g�l�F��H����V��L����u�l�u�k�u�m�F��I����W��_�E��d�e�d�e�u�}�W���O���F�_�D��e�e�d�e�g�l�G��H����W�d��U��g�h�u�e�f�l�F��I����V��_�E��d�d�d�y�]�}�W��Y���V��_�D��e�d�e�d�f�m�G��I����FǻN��L���k�w�e�d�f�m�G��H����V��_�E��d�w�u�u�w�k�B��Y����W��_�E��e�d�d�e�g�l�F��H���F�W�H���e�d�d�d�f�m�G��I����W��^�E��y�_�u�u�n�}�I���I����V��^�D��d�d�d�e�g�m�F���Y���P��S�W��d�d�e�e�g�l�F��I����W��^�W���u�u�c�l�j�}�G��H����V��_�E��d�e�d�e�g�l�[�ԜY����F�L�D��d�d�e�e�f�l�G��I����V��L����u�e�u�k�u�m�F��I����W��_�D��e�d�d�e�u�}�W���N���F�_�D��e�e�e�e�g�m�F��I����W�d��U��f�h�u�e�f�l�F��I����V��_�E��e�e�d�y�]�}�W��Y���V��_�D��d�e�d�e�f�l�F��I����FǻN��E���k�w�e�d�f�m�G��I����W��_�E��e�w�u�u�w�j�A��Y����W��_�E��e�d�e�d�f�l�F��I���F� ^�H���e�d�d�d�f�m�F��I����W��_�E��y�_�u�u�g�}�I���I����V��^�E��e�e�e�e�g�m�G���Y���Q��S�W��d�d�e�e�g�m�F��I����V��_�W���u�u�b�e�j�}�G��H����V��^�E��e�d�e�e�f�m�[�ԜY����F�L�D��d�d�e�d�g�l�F��I����V��L����u�d�u�k�u�m�F��I����V��^�E��d�d�e�d�u�}�W���N���F�_�D��e�e�e�e�f�m�G��H����V�d��U��a�h�u�e�f�l�F��I����V��^�E��e�e�d�y�]�}�W��Y���V��_�D��d�d�d�d�g�l�G��I����FǻN��D���k�w�e�d�f�m�G��I����W��_�E��d�w�u�u�w�j�@��Y����W��_�E��d�e�e�e�f�l�G��H���F� _�H���e�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�}�I���I����V��^�D��d�e�e�d�f�l�F���Y���Q��S�W��d�d�e�e�g�m�F��H����V��_�W���u�u�b�d�j�}�G��H����V��_�D��d�d�d�e�g�l�[�ԜY����F�L�D��d�d�e�d�f�l�F��I����W��L����u�g�u�k�u�m�F��I����W��^�E��e�e�e�d�u�}�W���N���F�_�D��e�e�d�e�f�l�F��H����V�d��U��`�h�u�e�f�l�F��I����W��^�E��e�d�d�y�]�}�W��Y���V��_�D��d�e�d�d�g�l�G��H����FǻN��G���k�w�e�d�f�m�G��H����V��_�D��e�w�u�u�w�j�O��Y����W��_�E��d�e�d�d�f�l�G��I���F� \�H���e�d�d�d�f�m�F��I����V��^�E��y�_�u�u�d�}�I���I����V��^�E��d�d�e�e�f�m�G���Y���Q��S�W��d�d�e�e�g�l�F��I����V��_�W���u�u�b�g�j�}�G��H����V��^�D��e�e�d�d�f�m�[�ԜY���� F�L�D��d�d�e�d�f�m�G��I����V��L����u�f�u�k�u�m�F��I����W��^�D��d�e�e�d�u�}�W���N���F�_�D��e�e�d�e�f�m�G��H����W�d��U��c�h�u�e�f�l�F��I����W��_�E��e�e�e�y�]�}�W��Y���V��_�D��d�d�d�e�f�l�G��H����FǻN��F���k�w�e�d�f�m�G��H����W��^�D��e�w�u�u�w�j�N��Y����W��_�E��d�e�e�e�g�l�F��I���F� Z�H���e�d�d�d�f�m�F��I����W��_�E��y�_�u�u�c�}�I���I����V��^�D��e�d�d�e�f�m�F���Y���Q��S�W��d�d�e�e�g�l�F��H����V��^�W���u�u�b�f�j�}�G��H����V��_�D��e�d�d�d�g�m�[�ԜY����F�L�D��d�d�e�e�g�m�G��I����W��L����u�a�u�k�u�m�F��I����V��_�D��e�d�e�d�u�}�W���N���F�_�D��e�d�e�e�f�l�F��I����W�d��U��b�h�u�e�f�l�F��I����W��_�E��d�e�d�y�]�}�W��Y���V��_�D��e�e�d�e�f�m�G��I����FǻN��A���k�w�e�d�f�m�G��I����V��_�E��e�w�u�u�w�j�G��Y����W��_�D��d�e�d�d�f�l�F��H���F� [�H���e�d�d�d�f�m�G��I����V��_�D��y�_�u�u�b�}�I���I����V��_�E��e�d�e�d�g�l�G���Y���Q��S�W��d�d�e�e�f�m�F��I����V��_�W���u�u�b�a�j�}�G��H����V��^�D��d�e�e�d�f�m�[�ԜY����F�L�D��d�d�e�e�f�m�F��H����W��L����u�`�u�k�u�m�F��I����V��_�D��d�e�e�e�u�}�W���N���F�_�D��e�d�e�e�g�m�F��I����W�d��U��m�h�u�e�f�l�F��I����W��_�E��e�d�d�y�]�}�W��Y���V��_�D��e�d�d�d�f�l�G��H����FǻN��C���k�w�e�d�f�m�G��I����W��_�D��e�w�u�u�w�j�F��Y����W��_�D��d�d�e�d�f�l�F��H���F� X�H���e�d�d�d�f�m�G��I����W��_�D��y�_�u�u�a�}�I���I����V��_�D��d�d�d�d�g�l�F���Y���Q��S�W��d�d�e�e�f�m�F��H����V��_�W���u�u�b�`�j�}�G��H����V��^�E��d�d�d�d�f�l�[�ԜY����F�L�D��d�d�e�e�g�m�F��H����W��L����u�c�u�k�u�m�F��I����W��_�E��e�e�e�d�u�}�W���N���F�_�D��e�d�d�e�g�m�G��I����W�d��U��l�h�u�e�f�l�F��I����W��^�E��e�e�d�y�]�}�W��Y���V��_�D��e�e�e�e�g�m�G��I����FǻN��B���k�w�e�d�f�m�G��H����W��^�D��e�w�u�u�w�j�E��Y����W��_�D��d�d�e�e�g�m�G��H���F� Y�H���e�d�d�d�f�m�G��H����V��_�E��y�_�u�u�`�}�I���I����V��_�E��e�e�e�d�f�m�F���Y���Q��S�W��d�d�e�e�f�l�F��H����W��^�W���u�u�b�c�j�}�G��H����V��_�E��e�e�d�d�g�m�[�ԜY����F�L�D��d�d�e�e�f�m�G��I����V��L����u�b�u�k�u�m�F��I����W��^�E��d�d�d�e�u�}�W���N���F�_�D��e�d�d�e�g�l�G��H����W�d��U��e�h�u�e�f�l�F��I����W��^�D��e�e�e�y�]�}�W��Y���V��_�D��e�d�e�e�g�m�G��H����FǻN��M���k�w�e�d�f�m�G��H����V��_�E��d�w�u�u�w�j�D��Y����W��_�D��d�d�d�e�f�m�F��H���F� V�H���e�d�d�d�f�m�G��H����V��^�D��y�_�u�u�o�}�I���I����V��_�D��e�e�e�e�g�l�G���Y���Q��S�W��d�d�e�e�f�m�G��I����V��^�W���u�u�b�b�j�}�G��H����V��^�E��e�d�e�d�g�m�[�ԜY����F�L�D��d�d�e�d�g�m�F��I����V��L����u�m�u�k�u�m�F��I����V��^�E��e�e�e�d�u�}�W���N���F�_�D��e�d�e�e�f�m�G��I����W�d��U��d�h�u�e�f�l�F��I����W��^�D��e�d�e�y�]�}�W��Y���V��_�D��d�e�e�d�g�m�F��H����FǻN��L���k�w�e�d�f�m�G��I����W��^�D��e�w�u�u�w�j�C��Y����W��_�D��d�e�e�e�g�l�G��H���F� W�H���e�d�d�d�f�m�F��H����V��^�D��y�_�u�u�n�}�I���I����V��_�E��d�e�e�d�g�l�F���Y���Q��S�W��d�d�e�e�f�m�G��H����V��_�W���u�u�b�m�j�}�G��H����V��_�D��e�e�e�e�f�l�[�ԜY����
F�L�D��d�d�e�d�f�m�F��I����W��L����u�e�u�k�u�m�F��I����V��^�E��d�e�e�d�u�}�W���A���F�_�D��e�d�e�e�f�l�G��H����V�d��U��g�h�u�e�f�l�F��I����V��^�E��d�e�d�y�]�}�W��Y���V��_�D��d�d�e�d�g�m�G��I����FǻN��E���k�w�e�d�f�m�G��I����V��^�D��d�w�u�u�w�e�B��Y����W��_�D��d�e�d�e�g�m�G��H���F�^�H���e�d�d�d�f�m�F��H����W��_�D��y�_�u�u�g�}�I���I����V��_�D��d�d�d�d�g�l�F���Y���^��S�W��d�d�e�e�f�l�G��H����V��_�W���u�u�m�l�j�}�G��H����V��^�D��d�d�e�e�f�l�[�ԜY����F�L�D��d�d�e�d�g�m�F��H����W��L����u�d�u�k�u�m�F��I����W��^�D��e�e�e�d�u�}�W���A���F�_�D��e�d�d�e�f�l�F��I����V�d��U��f�h�u�e�f�l�F��I����V��_�E��d�e�e�y�]�}�W��Y���V��_�D��d�e�e�d�f�l�F��H����FǻN��D���k�w�e�d�f�m�G��H����V��^�D��e�w�u�u�w�e�A��Y����W��_�D��d�e�d�d�g�l�F��I���F�_�H���e�d�d�d�f�m�F��H����W��^�E��y�_�u�u�f�}�I���I����V��_�E��d�d�d�e�g�l�F���Y���^��S�W��d�d�e�e�f�l�G��I����W��^�W���u�u�m�e�j�}�G��H����V��_�D��d�d�e�d�g�m�[�ԜY����F�L�D��d�d�e�d�f�l�G��I����V��L����u�g�u�k�u�m�F��I����W��^�D��e�e�d�d�u�}�W���A���F�_�D��e�d�d�e�f�m�F��I����V�d��U��a�h�u�e�f�l�F��I����V��_�E��d�d�d�y�]�}�W��Y���V��_�D��d�d�e�e�f�m�F��I����FǻN��G���k�w�e�d�f�m�G��H����W��^�D��d�w�u�u�w�e�@��Y����W��_�D��d�e�e�d�g�m�G��H���F�\�H���e�d�d�d�f�m�F��H����W��_�D��y�_�u�u�e�}�I���I����V��^�E��e�d�d�d�f�l�F���Y���^��S�W��d�d�e�e�g�m�G��H����W��_�W���u�u�m�d�j�}�G��H����W��^�D��e�d�e�e�g�l�[�ԜY����F�L�D��d�d�d�e�g�l�G��H����V��L����u�f�u�k�u�m�F��I����V��_�D��d�e�d�d�u�}�W���A���F�_�D��e�e�e�e�f�l�G��H����W�d��U��`�h�u�e�f�l�F��H����V��_�E��e�d�d�y�]�}�W��Y���V��_�D��e�e�e�e�f�m�F��I����FǻN��F���k�w�e�d�f�m�G��I����V��_�D��d�w�u�u�w�e�O��Y����W��_�E��d�e�d�e�f�m�G��I���F�]�H���e�d�d�d�f�l�G��H����V��^�E��y�_�u�u�c�}�I���I����V��^�D��e�d�e�d�g�m�F���Y���^��S�W��d�d�e�e�g�m�G��I����V��_�W���u�u�m�g�j�}�G��H����W��_�D��d�d�d�e�g�m�[�ԜY���� F�L�D��d�d�d�e�f�l�F��H����W��L����u�a�u�k�u�m�F��I����V��_�E��e�d�e�d�u�}�W���A���F�_�D��e�e�e�d�g�m�F��H����V�d��U��c�h�u�e�f�l�F��H����V��^�E��d�d�d�y�]�}�W��Y���V��_�D��e�d�e�d�g�l�G��I����FǻN��A���k�w�e�d�f�m�G��I����W��_�E��e�w�u�u�w�e�N��Y����W��_�E��d�d�e�d�f�l�G��I���F�[�H���e�d�d�d�f�l�G��H����V��^�D��y�_�u�u�b�}�I���I����V��^�E��d�e�e�d�f�m�F���Y���^��S�W��d�d�e�e�g�l�G��H����V��_�W���u�u�m�f�j�}�G��H����W��^�E��e�d�d�d�g�l�[�ԜY����F�L�D��d�d�d�e�g�l�F��H����V��L����u�`�u�k�u�m�F��I����W��_�E��e�e�d�e�u�}�W���A���F�_�D��e�e�d�d�g�l�G��I����W�d��U��b�h�u�e�f�l�F��H����V��^�E��d�e�d�y�]�}�W��Y���V��_�D��e�e�e�d�g�m�F��I����FǻN��@���k�w�e�d�f�m�G��H����V��_�E��d�w�u�u�w�e�G��Y����W��_�E��d�d�d�e�g�l�G��H���F�X�H���e�d�d�d�f�l�G��I����V��_�E��y�_�u�u�a�}�I���I����V��^�D��d�d�d�d�f�l�F���Y���^��S�W��d�d�e�e�g�l�G��H����V��^�W���u�u�m�a�j�}�G��H����W��_�E��d�d�e�d�g�m�[�ԜY����F�L�D��d�d�d�e�f�l�F��H����W��L����u�c�u�k�u�m�F��I����W��_�D��e�e�d�d�u�}�W���A���F�_�D��e�e�d�d�g�l�F��I����W�d��U��m�h�u�e�f�l�F��H����V��_�D��e�d�d�y�]�}�W��Y���V��_�D��e�d�e�d�f�m�F��I����FǻN��B���k�w�e�d�f�m�G��H����V��^�D��e�w�u�u�w�e�F��Y����W��_�E��d�d�d�e�f�m�G��H���F�Y�H���e�d�d�d�f�l�F��I����W��^�D��y�_�u�u�`�}�I���I����V��^�E��d�d�d�d�g�l�G���Y���^��S�W��d�d�e�e�g�m�G��I����V��^�W���u�u�m�`�j�}�G��H����W��^�E��e�d�e�e�g�l�[�ԜY����F�L�D��d�d�d�d�g�l�G��I����W��L����u�b�u�k�u�m�F��I����V��_�D��e�d�e�d�u�}�W���A���F�_�D��e�e�e�d�g�m�F��H����W�d��U��l�h�u�e�f�l�F��H����V��^�D��d�d�d�y�]�}�W��Y���V��_�D��d�e�d�e�g�l�F��I����FǻN��M���k�w�e�d�f�m�G��I����W��^�D��e�w�u�u�w�e�E��Y����W��_�E��d�d�e�d�f�m�F��H���F�V�H���e�d�d�d�f�l�F��I����V��^�D��y�_�u�u�o�}�I���I����V��^�D��e�e�e�e�f�l�F���Y���^��S�W��d�d�e�e�g�m�G��H����W��_�W���u�u�m�c�j�}�G��H����W��_�E��e�d�e�d�g�l�[�ԜY����F�L�D��d�d�d�d�f�l�G��H����W��L����u�m�u�k�u�m�F��I����V��^�E��e�e�e�e�u�}�W���A���F�_�D��e�e�e�d�g�l�G��H����W�d��U��e�h�u�e�f�l�F��H����V��^�E��d�d�d�y�]�}�W��Y���V��_�D��d�d�d�e�g�m�G��H����FǻN��L���k�w�e�d�f�m�G��I����W��_�D��d�w�u�u�w�e�D��Y����W��_�E��d�d�e�d�g�l�F��H���F�W�H���e�d�d�d�f�l�F��I����W��_�E��y�_�u�u�n�}�I���I����V��^�E��e�d�e�e�f�l�F���Y���^��S�W��d�d�e�e�g�l�G��H����W��_�W���u�u�m�b�j�}�G��H����W��^�E��d�e�e�e�f�l�[�ԜY����F�L�D��d�d�d�d�g�l�G��H����W��L����u�l�u�k�u�m�F��I����W��^�D��d�e�e�d�u�}�W���@���F�_�D��e�e�d�d�g�l�G��I����W�d��U��d�h�u�e�f�l�F��H����V��_�D��e�e�e�y�]�}�W��Y���V��_�D��d�e�d�e�f�m�F��H����FǻN��E���k�w�e�d�f�m�G��H����V��_�D��e�w�u�u�w�d�C��Y����W��_�E��d�d�d�d�f�m�F��I���F�^�H���e�d�d�d�f�l�F��I����W��^�E��y�_�u�u�g�}�I���I����V��^�D��e�e�e�d�g�m�F���Y���_��S�W��d�d�e�e�g�l�G��I����V��^�W���u�u�l�m�j�}�G��H����W��_�E��d�e�d�e�g�l�[�ԜY����
F�L�D��d�d�d�d�f�l�F��H����V��L����u�d�u�k�u�m�F��I����W��^�E��d�e�e�e�u�}�W���@���F�_�D��e�e�d�d�f�m�G��I����V�d��U��g�h�u�e�f�l�F��H����V��^�D��d�e�e�y�]�}�W��Y���V��_�D��d�d�d�d�g�m�G��I����FǻN��D���k�w�e�d�f�m�G��H����V��_�D��e�w�u�u�w�d�B��Y����W��_�E��d�d�d�d�g�l�F��H���F�_�H���e�d�d�d�f�l�G��I����W��^�E��y�_�u�u�f�}�I���I����V��_�E��e�d�e�e�g�m�G���Y���_��S�W��d�d�e�e�f�m�G��I����W��^�W���u�u�l�l�j�}�G��H����W��^�E��e�d�e�d�f�l�[�ԜY����F�L�D��d�d�d�e�g�l�F��H����W��L����u�g�u�k�u�m�F��I����V��^�D��d�d�e�e�u�}�W���@���F�_�D��e�d�e�d�f�m�G��I����V�d��U��f�h�u�e�f�l�F��H����V��_�E��e�d�d�y�]�}�W��Y���V��_�D��e�e�d�d�g�l�G��H����FǻN��G���k�w�e�d�f�m�G��I����W��^�E��d�w�u�u�w�d�A��Y����W��_�D��e�e�e�d�f�m�F��I���F�\�H���e�d�d�d�f�l�G��I����V��^�E��y�_�u�u�e�}�I���I����V��_�D��d�e�d�d�f�l�F���Y���_��S�W��d�d�e�e�f�m�G��H����V��_�W���u�u�l�e�j�}�G��H����W��_�D��e�e�e�e�f�l�[�ԜY����F�L�D��d�d�d�e�f�l�F��I����V��L����u�f�u�k�u�m�F��I����V��^�E��e�e�d�e�u�}�W���@���F�_�D��e�d�e�d�f�m�F��H����V�d��U��a�h�u�e�f�l�F��H����V��_�E��e�e�e�y�]�}�W��Y���V��_�D��e�d�d�d�f�m�F��I����FǻN��F���k�w�e�d�f�m�G��I����W��^�D��e�w�u�u�w�d�@��Y����W��_�D��e�e�e�e�f�m�F��I���F�]�H���e�d�d�d�f�l�G��I����W��^�E��y�_�u�u�d�}�I���I����V��_�E��d�d�e�d�g�l�G���Y���_��S�W��d�d�e�e�f�l�G��H����W��_�W���u�u�l�d�j�}�G��H����W��^�D��d�d�d�d�f�m�[�ԜY����F�L�D��d�d�d�e�g�l�F��H����V��L����u�a�u�k�u�m�F��I����W��^�E��d�d�d�e�u�}�W���@���F�_�D��e�d�d�d�f�l�F��H����V�d��U��`�h�u�e�f�l�F��H����W��^�D��e�d�d�y�]�}�W��Y���V��_�D��e�e�d�d�g�l�F��H����FǻN��A���k�w�e�d�f�m�G��H����V��_�D��d�w�u�u�w�d�O��Y����W��_�D��e�e�d�e�g�l�G��I���F�Z�H���e�d�d�d�f�l�G��I����W��_�E��y�_�u�u�b�}�I���I����V��_�D��d�d�d�d�g�l�G���Y���_��S�W��d�d�e�e�f�l�G��H����W��_�W���u�u�l�g�j�}�G��H����W��_�D��d�e�d�e�g�l�[�ԜY���� F�L�D��d�d�d�e�f�l�F��H����V��L����u�`�u�k�u�m�F��I����W��^�D��d�d�e�d�u�}�W���@���F�_�D��e�d�d�d�f�l�G��I����W�d��U��c�h�u�e�f�l�F��H����W��_�E��e�d�e�y�]�}�W��Y���V��_�D��e�d�d�d�g�l�G��I����FǻN��@���k�w�e�d�f�m�G��H����V��^�E��d�w�u�u�w�d�N��Y����W��_�D��e�e�d�d�f�l�G��H���F�X�H���e�d�d�d�f�l�F��I����V��_�E��y�_�u�u�a�}�I���I����V��_�E��d�e�d�e�g�l�F���Y���_��S�W��d�d�e�e�f�m�G��I����W��^�W���u�u�l�f�j�}�G��H����W��^�D��e�e�d�d�g�l�[�ԜY����F�L�D��d�d�d�d�g�l�F��H����V��L����u�c�u�k�u�m�F��I����V��^�D��d�e�e�e�u�}�W���@���F�_�D��e�d�e�d�f�l�F��H����V�d��U��b�h�u�e�f�l�F��H����W��_�E��e�d�e�y�]�}�W��Y���V��_�D��d�e�d�d�f�l�G��H����FǻN��C���k�w�e�d�f�m�G��I����V��_�D��e�w�u�u�w�d�G��Y����W��_�D��e�e�d�e�g�l�G��I���F�Y�H���e�d�d�d�f�l�F��I����W��^�D��y�_�u�u�`�}�I���I����V��_�D��d�e�d�e�f�l�F���Y���_��S�W��d�d�e�e�f�m�G��I����V��_�W���u�u�l�a�j�}�G��H����W��_�D��d�e�e�e�g�l�[�ԜY����F�L�D��d�d�d�d�f�m�G��H����V��L����u�b�u�k�u�m�F��I����V��^�E��d�d�e�e�u�}�W���@���F�_�D��e�d�e�d�f�m�G��H����W�d��U��m�h�u�e�f�l�F��H����W��_�D��e�d�d�y�]�}�W��Y���V��_�D��d�d�d�d�f�m�F��I����FǻN��M���k�w�e�d�f�m�G��I����V��^�D��d�w�u�u�w�d�F��Y����W��_�D��e�e�d�e�f�l�F��H���F�V�H���e�d�d�d�f�l�F��I����W��_�D��y�_�u�u�o�}�I���I����V��_�E��d�d�e�d�f�m�G���Y���_��S�W��d�d�e�e�f�l�G��I����V��_�W���u�u�l�`�j�}�G��H����W��^�D��d�e�d�e�g�l�[�ԜY����F�L�D��d�d�d�d�g�m�G��I����V��L����u�m�u�k�u�m�F��I����W��^�E��d�e�e�d�u�}�W���@���F�_�D��e�d�d�d�f�m�G��I����W�d��U��l�h�u�e�f�l�F��H����W��^�D��d�d�d�y�]�}�W��Y���V��_�D��d�e�d�d�f�l�F��H����FǻN��L���k�w�e�d�f�m�G��H����V��^�E��e�w�u�u�w�d�E��Y����W��_�D��e�e�d�d�f�l�G��I���F�W�H���e�d�d�d�f�l�F��I����W��_�D��y�_�u�u�n�}�I���I����V��_�D��d�d�d�d�g�l�F���Y���_��S�W��d�d�e�e�f�l�G��I����W��_�W���u�u�l�c�j�}�G��H����W��_�D��d�d�d�e�g�l�[�ԜY����F�L�D��d�d�d�d�f�m�G��H����W��L����u�l�u�k�u�m�F��I����W��^�E��e�d�e�e�u�}�W���@���F�_�D��e�d�d�d�f�m�G��H����V�d��U��e�u�k�w�g�l�F��I����W��_�D��d�d�d�w�w�}�W��I���D��_�D��d�d�d�d�g�m�G��I����D�=N��U��g�h�u�e�f�l�F��H����W��_�D��e�d�d�y�]�}�W��J���V��_�E��e�e�e�e�f�l�G��H����J�N��D��u�k�w�e�f�l�G��I����W��_�D��e�e�w�u�w�}�F��Y���V��_�D��e�e�e�d�f�l�G��H����FǻN��E��h�u�e�d�f�l�F��I����W��^�D��d�d�y�_�w�}�G��D���W��_�D��e�e�d�d�g�m�G��H���l�N�E���k�w�e�d�f�m�F��I����V��_�E��d�w�u�u�w�l�G���G����W��^�E��e�e�d�e�g�l�F��H���9F�_�E��u�e�d�d�f�l�G��I����V��^�D��d�y�_�u�w�m�F��Y����W��_�E��d�e�d�e�g�l�G��I���F�^�U��w�e�d�d�g�l�G��H����V��_�D��w�u�u�u�f�l�W���[����W��_�E��d�d�d�d�f�m�F��[��ƹF�_�H���e�d�d�d�f�m�G��I����W��^�E��y�_�u�u�g�h�J���I����W��^�E��d�e�d�e�f�l�F��U���F��X��K���e�d�d�e�f�m�G��H����W��_�E���u�u�u�d�f�}�I���I����V��^�D��d�d�e�d�g�m�G���Y���W��N��U��d�d�d�d�g�m�F��I����V��^�D���_�u�u�e�n�`�W��H����W��^�D��e�d�e�d�g�m�F��s���V��S�W��d�d�e�d�g�m�F��H����W��_�W���u�u�d�g�w�c�U��H����W��^�E��e�d�d�d�f�l�U���Y���T��
P��E��d�d�d�e�g�l�F��I����W��^�Y�ߊu�u�e�f�j�}�G��H����V��_�D��e�e�e�e�f�m�[�ԜY����R�	N��E��d�e�d�e�g�l�F��H����W��_��U���u�d�g�u�i��G��H����V��^�E��e�d�e�e�g��W���Y����F�L�D��d�d�e�e�g�m�G��H����V��L����u�e�b�h�w�m�F��H����V��^�D��e�d�d�d�g�q�}���Y����[�^�D��e�d�e�d�g�m�G��I����V��B��U���d�g�u�k�u�m�F��I����W��_�E��e�d�e�e�u�}�W���H����X�^�D��d�e�e�e�g�m�G��H����W��NךU���e�d�h�u�g�l�F��H����V��_�E��d�d�e�e�{�W�W���I���F�_�D��d�e�d�d�f�m�G��H����V�d��U��f�u�k�w�g�l�F��H����W��_�E��d�d�e�w�w�}�W��J���D��_�D��e�e�e�d�f�l�F��I����D�=N��U��`�h�u�e�f�l�F��I����W��_�D��d�d�d�y�]�}�W��O���V��_�E��e�d�e�e�f�m�F��H����J�N��D��u�k�w�e�f�l�G��I����W��^�E��d�d�w�u�w�}�F��Y���V��_�D��e�d�e�d�f�m�F��I����FǻN��E��h�u�e�d�f�l�F��I����W��_�D��d�e�y�_�w�}�G��D���W��_�D��d�e�d�d�f�l�G��I���l�N�A���k�w�e�d�f�m�F��H����V��_�D��d�w�u�u�w�l�C���G����W��^�E��d�e�d�e�g�l�G��H���9F�_�F��u�e�d�d�f�l�G��H����V��^�D��d�y�_�u�w�m�C��Y����W��_�E��d�e�e�d�g�l�G��I���F�^�U��w�e�d�d�g�l�G��H����W��^�D��w�u�u�u�f�i�W���[����W��_�E��d�d�d�d�f�l�G��[��ƹF�Z�H���e�d�d�d�f�m�F��I����V��_�E��y�_�u�u�g�e�J���I����W��^�E��d�e�d�d�f�l�F��U���F��W��K���e�d�d�e�f�m�G��H����W��_�D���u�u�u�d�b�}�I���I����V��^�E��d�e�d�d�f�l�G���Y���W��N��U��d�d�d�d�g�l�G��I����V��_�D���_�u�u�e�e�`�W��H����W��_�D��e�e�e�d�f�l�F��s���V��S�W��d�d�e�d�g�m�F��I����V��^�W���u�u�d�`�w�c�U��H����W��^�E��d�e�d�d�f�m�U���Y���S��
P��E��d�d�d�e�f�m�F��H����V��_�Y�ߊu�u�e�c�j�}�G��H����V��^�E��e�d�d�d�g�l�[�ԜY����Q�	N��E��d�e�d�e�g�l�F��H����V��_��U���u�d�`�u�i��G��H����V��^�E��e�d�d�e�g��W���Y����
F�L�D��d�d�e�d�f�m�G��H����V��L����u�e�e�h�w�m�F��H����W��^�D��e�e�d�e�g�q�}���Y����[�^�D��e�d�e�e�g�m�G��I����V��B��U���d�c�u�k�u�m�F��I����V��_�D��e�d�e�d�u�}�W���H����X�^�D��d�e�d�d�f�l�F��H����V��NךU���e�a�h�u�g�l�F��H����W��_�E��e�e�d�e�{�W�W���I���F�_�D��d�e�e�d�f�l�G��H����V�d��U��c�u�k�w�g�l�F��H����W��^�D��d�e�e�w�w�}�W��O���D��_�D��e�d�d�d�f�m�G��I����D�=N��U��m�h�u�e�f�l�F��I����W��^�D��e�d�e�y�]�}�W��@���V��_�E��e�d�e�e�f�m�F��I����J�N��D��u�k�w�e�f�l�G��I����V��_�E��e�e�w�u�w�}�F��Y���V��_�D��d�e�e�d�f�m�G��I����FǻN��E��h�u�e�d�f�l�F��H����V��_�E��e�d�y�_�w�}�G��D���W��_�D��d�e�d�e�g�l�G��H���l�N�B���k�w�e�d�f�m�F��H����W��_�D��d�w�u�u�w�l�@���G����W��^�E��e�e�d�e�g�l�F��H���9F�_�C��u�e�d�d�f�l�G��I����V��_�E��e�y�_�u�w�m�@��Y����W��_�E��d�e�e�e�f�l�F��H���F�^�U��w�e�d�d�g�l�G��H����W��_�D��w�u�u�u�f�j�W���[����W��_�D��d�e�d�e�f�l�G��[��ƹF�V�H���e�d�d�d�f�m�F��I����W��_�E��y�_�u�u�g�l�J���I����W��^�D��e�d�e�d�f�m�F��U���F��\��K���e�d�d�e�f�m�F��H����W��^�D���u�u�u�d�o�}�I���I����V��^�D��e�e�e�d�f�l�G���Y���W��N��U��d�d�d�d�g�l�F��I����W��_�E���_�u�u�e�b�`�W��H����W��_�E��d�e�d�d�g�l�F��s���V��S�W��d�d�e�d�g�l�F��H����W��_�W���u�u�d�m�w�c�U��H����W��_�E��d�e�d�e�g�m�U���Y���^��
P��E��d�d�d�e�f�l�G��H����V��_�Y�ߊu�u�e�l�j�}�G��H����V��_�E��e�d�e�d�f�l�[�ԜY����
V�	N��E��d�e�d�e�f�l�F��H����V��^��U���u�d�l�u�i��G��H����W��^�E��e�d�e�d�g��W���Y����F�L�D��d�d�e�e�g�m�F��H����W��L����u�e�f�h�w�m�F��H����V��^�E��d�d�d�d�f�q�}���Y����[�^�D��e�d�d�e�g�m�G��H����W��B��U���d�l�u�k�u�m�F��I����V��^�D��e�e�e�e�u�}�W���H����X�^�D��d�e�e�e�f�l�F��I����W��NךU���e�b�h�u�g�l�F��H����V��^�E��e�e�d�d�{�W�W���I���F�_�D��d�d�e�d�f�m�F��H����V�d��U��l�u�k�w�g�l�F��H����W��_�E��e�d�e�w�w�}�W��I���D��_�D��e�e�e�d�f�m�F��H����D�=N��U��d�h�u�e�f�l�F��I����W��^�E��e�d�d�y�]�}�W��K���V��_�E��d�e�d�d�f�l�G��H����J�N��D��u�k�w�e�f�l�G��H����V��_�E��e�e�w�u�w�}�F��Y���V��_�D��e�d�e�e�f�l�G��H����FǻN��D���h�u�e�d�f�l�F��I����V��_�D��d�e�y�_�w�}�F��D���W��_�D��e�e�e�d�f�l�G��H���l�N�E���k�w�e�d�f�m�F��I����V��_�D��e�w�u�u�w�l�G���G����W��^�E��d�e�e�e�g�m�G��I���9F�_�L��u�e�d�d�f�l�G��H����W��^�D��d�y�_�u�w�l�G��Y����W��_�D��d�d�e�d�g�l�F��H���F�_�U��w�e�d�d�g�l�F��H����V��^�E��w�u�u�u�f�l�W���[����W��_�E��d�e�d�e�g�l�G��[��ƹF�_�H���e�d�d�d�f�m�G��H����W��_�E��y�_�u�u�f�i�J���I����W��^�D��e�e�e�d�f�m�G��U���F��[��K���e�d�d�e�f�l�F��H����W��^�E���u�u�u�d�f�}�I���I����V��_�E��d�d�d�e�f�m�G���Y���W�� N��U��d�d�d�d�g�m�G��H����V��_�D���_�u�u�d�o�`�W��H����W��^�E��d�e�e�d�f�l�F��s���W��S�W��d�d�e�d�f�l�F��I����V��_�W���u�u�d�g�w�c�U��H����W��_�E��e�d�e�e�g�m�U���Y���T��
P��E��d�d�d�e�g�m�G��I����W��_�Y�ߊu�u�d�g�j�}�G��H����V��^�E��e�d�e�e�f�m�[�ԜY����U�	N��E��d�e�d�d�f�l�G��H����W��^��U���u�d�g�u�i��G��H����W��_�D��e�d�d�d�g��W���Y����F�L�D��d�d�e�e�f�m�G��H����V��L����u�d�c�h�w�m�F��H����V��^�E��e�d�e�d�f�q�}���Y����[�^�D��e�d�d�d�g�l�F��H����W��B��U���d�g�u�k�u�m�F��I����W��^�E��d�e�d�e�u�}�W���H����X�^�D��d�e�e�d�f�m�G��I����W��NךU���d�e�h�u�g�l�F��H����W��_�D��d�d�e�e�{�W�W���H���F�_�D��d�d�d�d�g�m�F��H����W�d��U��f�u�k�w�g�l�F��H����W��_�D��e�e�d�w�w�}�W��J���D��_�D��e�e�d�d�g�m�F��H����D�=N��U��a�h�u�e�f�l�F��I����W��^�D��e�e�d�y�]�}�W��L���V��_�E��d�d�d�d�g�m�G��H����J�N��D��u�k�w�e�f�l�G��H����V��^�E��d�d�w�u�w�}�F��Y���V��_�D��d�e�e�d�f�m�F��H����FǻN��D��h�u�e�d�f�l�F��H����W��_�E��e�d�y�_�w�}�F��D���W��_�D��e�e�e�d�g�l�G��I���l�N�A���k�w�e�d�f�m�F��I����V��^�D��d�w�u�u�w�l�C���G����W��^�E��e�d�d�e�g�m�F��I���9F�_�G��u�e�d�d�f�l�G��I����V��_�D��e�y�_�u�w�l�D��Y����W��_�D��d�d�e�d�f�m�F��H���F�_�U��w�e�d�d�g�l�F��H����W��^�D��w�u�u�u�f�i�W���[����W��_�D��d�d�d�d�g�l�F��[��ƹF�Z�H���e�d�d�d�f�m�F��H����W��_�D��y�_�u�u�f�j�J���I����W��^�E��e�e�d�d�g�l�G��U���F��V��K���e�d�d�e�f�l�G��I����V��^�E���u�u�u�d�c�}�I���I����V��_�D��d�e�e�e�f�m�G���Y���W��N��U��d�d�d�d�g�l�F��I����W��_�D���_�u�u�d�f�`�W��H����W��_�E��d�e�d�e�g�l�F��s���W��S�W��d�d�e�d�f�m�G��I����V��^�W���u�u�d�`�w�c�U��H����W��^�E��e�e�d�d�g�m�U���Y���S��
P��E��d�d�d�e�f�l�G��I����V��^�Y�ߊu�u�d�`�j�}�G��H����V��_�D��e�e�d�e�g�m�[�ԜY����P�	N��E��d�e�d�d�g�l�G��H����W��_��U���u�d�`�u�i��G��H����W��_�E��d�d�e�d�g��W���Y����F�L�D��d�d�e�d�f�l�F��I����W��L����u�d�l�h�w�m�F��H����W��^�E��e�d�e�e�g�q�}���Y����[�^�D��e�d�d�d�g�l�F��H����V��B��U���d�c�u�k�u�m�F��I����W��^�E��e�e�d�d�u�}�W���H����X�^�D��d�e�d�e�f�l�F��I����V��NךU���d�f�h�u�g�l�F��H����V��^�E��d�d�d�e�{�W�W���H���F�_�D��d�d�d�d�g�m�G��I����V�d��U��c�u�k�w�g�l�F��H����W��_�D��e�e�e�w�w�}�W��O���D��_�D��e�d�e�e�f�m�F��I����D�=N��U��b�h�u�e�f�l�F��I����W��^�D��e�e�e�y�]�}�W��A���V��_�E��d�d�d�e�f�l�G��H����J�N��D��u�k�w�e�f�l�G��H����W��^�D��e�d�w�u�w�}�F��Y���V��_�D��d�d�e�e�f�m�G��I����FǻN��D��h�u�e�d�f�l�F��H����V��_�D��e�d�y�_�w�}�F��D���W��_�D��d�e�d�d�g�l�G��I���l�N�B���k�w�e�d�f�m�F��H����V��^�D��d�w�u�u�w�l�@���G����W��^�E��d�d�e�d�f�m�F��H���9F�_�@��u�e�d�d�f�l�G��H����W��^�E��e�y�_�u�w�l�A��Y����W��_�D��d�e�e�e�g�m�G��H���F�_�U��w�e�d�d�g�l�F��H����W��_�E��w�u�u�u�f�j�W���[����W��_�D��d�e�e�d�g�m�F��[��ƹF�Y�H���e�d�d�d�f�m�F��H����V��^�D��y�_�u�u�f�m�J���I����W��^�D��d�d�d�d�g�m�F��U���F��_��K���e�d�d�e�f�m�G��I����V��^�E���u�u�u�d�o�}�I���I����V��^�E��d�e�d�d�f�m�F���Y���W��N��U��d�d�d�d�f�m�G��H����V��^�E���_�u�u�d�c�`�W��H����W��^�E��d�e�e�d�g�l�F��s���W��S�W��d�d�e�d�g�m�G��H����W��^�W���u�u�d�m�w�c�U��H����W��^�D��d�e�d�d�g�l�U���Y���^��
P��E��d�d�d�d�g�m�G��H����V��^�Y�ߊu�u�d�m�j�}�G��H����W��^�D��d�e�d�e�f�m�[�ԜY����_�	N��E��d�e�d�e�g�l�F��H����W��^��U���u�d�l�u�i��G��H����V��_�D��e�e�d�e�g��W���Y����F�L�D��d�d�d�e�g�l�G��H����W��L����u�d�g�h�w�m�F��H����V��_�D��d�d�e�e�g�q�}���Y����[�^�D��e�d�e�e�g�m�G��I����W��B��U���d�l�u�k�u�m�F��I����V��_�E��d�e�d�d�u�}�W���H����X�^�D��d�d�e�d�f�m�G��H����V��NךU���d�c�h�u�g�l�F��H����W��_�D��d�e�d�e�{�W�W���H���F�_�D��d�e�e�e�f�l�F��H����W�d��U��l�u�k�w�g�l�F��H����W��^�E��d�e�d�w�w�}�W��@���D��_�D��d�e�d�e�f�m�F��H����D�=N��U��e�h�u�e�f�l�F��H����V��^�D��d�e�e�y�]�}�W��H���V��_�E��e�e�d�e�f�m�F��I����J�N��D��u�k�w�e�f�l�G��I����V��_�E��d�e�w�u�w�}�F��Y���V��_�D��e�d�d�d�f�l�G��H����FǻN��G��h�u�e�d�f�l�F��I����V��^�E��d�e�y�_�w�}�E��D���W��_�D��d�e�d�e�f�l�G��H���l�N�E���k�w�e�d�f�m�F��H����W��^�E��d�w�u�u�w�l�G���G����W��^�D��e�d�e�d�f�m�G��I���9F�_�M��u�e�d�d�f�l�F��I����W��_�D��e�y�_�u�w�o�N��Y����W��_�E��e�d�d�e�g�l�F��H���F�\�U��w�e�d�d�g�l�G��H����W��_�D��w�u�u�u�f�l�W���[����W��_�E��e�e�e�d�f�m�F��[��ƹF�_�H���e�d�d�d�f�l�G��I����W��^�E��y�_�u�u�e�n�J���I����W��_�D��e�e�d�e�g�l�G��U���F��Z��K���e�d�d�e�f�m�F��H����W��^�E���u�u�u�d�f�}�I���I����V��^�D��e�e�d�d�g�l�F���Y���W��N��U��d�d�d�d�f�m�F��H����V��^�D���_�u�u�g�`�`�W��H����W��^�E��e�e�e�d�f�m�G��s���T��S�W��d�d�e�d�g�l�G��I����V��_�W���u�u�d�d�w�c�U��H����W��_�D��d�d�e�e�f�m�U���Y���T��
P��E��d�d�d�d�g�l�F��I����W��_�Y�ߊu�u�g�d�j�}�G��H����W��_�E��e�d�d�d�f�l�[�ԜY����T�	N��E��d�e�d�e�f�l�F��I����W��_��U���u�d�g�u�i��G��H����V��_�D��e�d�e�d�g��W���Y����F�L�D��d�d�d�e�f�l�G��H����W��L����u�g�`�h�w�m�F��H����V��_�E��d�e�d�e�f�q�}���Y����[�^�D��e�d�e�d�f�l�F��I����V��B��U���d�g�u�k�u�m�F��I����V��^�E��d�e�e�e�u�}�W���H����X�^�D��d�d�d�e�g�m�F��H����V��NךU���g�l�h�u�g�l�F��H����V��_�E��d�e�d�e�{�W�W���K���F�_�D��d�e�e�e�g�m�F��I����V�d��U��f�u�k�w�g�l�F��H����V��_�D��d�e�e�w�w�}�W��J���D��_�D��d�d�e�e�g�m�G��H����D�=N��U��f�h�u�e�f�l�F��H����V��_�D��d�e�e�y�]�}�W��M���V��_�E��e�e�d�d�f�m�G��H����J�N��D��u�k�w�e�f�l�G��I����V��_�D��e�e�w�u�w�}�F��Y���V��_�D��d�e�d�d�g�l�F��H����FǻN��G��h�u�e�d�f�l�F��H����W��^�D��d�e�y�_�w�}�E��D���W��_�D��e�e�e�e�f�l�G��H���l�N�F���k�w�e�d�f�m�F��I����W��_�E��e�w�u�u�w�l�C���G����W��^�D��d�e�d�e�f�l�G��I���9F�_�D��u�e�d�d�f�l�F��H����V��^�D��e�y�_�u�w�o�E��Y����W��_�E��e�e�d�d�f�l�F��H���F�\�U��w�e�d�d�g�l�G��I����W��^�D��w�u�u�u�f�i�W���[����W��_�D��e�e�d�e�g�l�G��[��ƹF�Z�H���e�d�d�d�f�l�F��I����V��^�D��y�_�u�u�e�k�J���I����W��_�E��d�d�e�e�f�l�G��U���F��Y��K���e�d�d�e�f�m�G��I����W��_�E���u�u�u�d�c�}�I���I����V��^�D��e�d�d�d�f�l�F���Y���W��N��U��d�d�d�d�f�l�F��H����V��_�E���_�u�u�g�g�`�W��H����W��_�E��e�d�e�d�f�m�F��s���T��S�W��d�d�e�d�g�l�G��H����V��^�W���u�u�d�`�w�c�U��H����W��_�E��d�d�e�d�g�m�U���Y���S��
P��E��d�d�d�d�f�m�F��H����W��^�Y�ߊu�u�g�a�j�}�G��H����W��^�D��d�d�d�e�f�l�[�ԜY����S�	N��E��d�e�d�e�f�l�G��I����W��^��U���u�d�`�u�i��G��H����V��_�D��e�e�d�e�f��W���Y����F�L�D��d�d�d�d�g�m�G��I����W��L����u�g�m�h�w�m�F��H����W��_�E��d�d�d�d�g�q�}���Y����[�^�D��e�d�e�d�f�m�F��H����W��B��U���d�c�u�k�u�m�F��I����W��_�E��d�e�e�e�u�}�W���H����X�^�D��d�d�d�d�g�m�F��I����W��NךU���g�g�h�u�g�l�F��H����W��_�E��e�e�e�d�{�W�W���K���F�_�D��d�e�d�e�f�m�F��H����V�d��U��c�u�k�w�g�l�F��H����V��_�E��d�d�e�w�w�}�W��O���D��_�D��d�d�d�d�g�m�G��H����D�=N��U��c�h�u�e�f�l�F��H����W��_�D��e�d�d�y�]�}�W��N���V��_�E��e�d�d�e�f�m�F��H����J�N��D��u�k�w�e�f�l�G��I����W��_�E��d�e�w�u�w�}�F��Y���V��_�D��d�d�e�d�g�l�F��H����FǻN��G��h�u�e�d�f�l�F��H����V��_�E��e�e�y�_�w�}�E��D���W��_�D��d�d�d�e�g�l�G��I���l�N�B���k�w�e�d�f�m�F��H����W��_�D��d�w�u�u�w�l�@���G����W��^�D��e�e�d�e�g�m�F��I���9F�_�A��u�e�d�d�f�l�F��I����V��_�E��d�y�_�u�w�o�B��Y����W��_�D��e�d�d�d�f�m�G��I���F�\�U��w�e�d�d�g�l�F��I����V��^�E��w�u�u�u�f�j�W���[����W��_�E��d�e�e�e�f�l�G��[��ƹF�Y�H���e�d�d�d�f�l�G��I����W��_�D��y�_�u�u�e�d�J���I����W��_�E��e�e�d�e�g�l�F��U���F��^��K���e�d�d�e�f�l�G��H����V��^�D���u�u�u�d�o�}�I���I����V��_�E��e�e�d�e�f�l�G���Y���W��N��U��d�d�d�d�f�m�G��H����W��_�E���_�u�u�g�d�`�W��H����W��^�D��d�d�d�d�f�l�F��s���T��S�W��d�d�e�d�f�m�G��I����V��^�W���u�u�d�m�w�c�U��H����W��^�E��d�e�e�d�g�l�U���Y���^��
P��E��d�d�d�d�g�l�G��I����W��_�Y�ߊu�u�g�b�j�}�G��H����W��_�E��e�d�e�e�g�m�[�ԜY����^�	N��E��d�e�d�d�g�m�G��H����V��_��U���u�d�m�u�i��G��H����W��^�D��e�d�e�e�g��W���Y����F�L�D��d�d�d�e�f�m�G��I����V��L����u�g�d�h�w�m�F��H����V��^�E��d�d�d�d�g�q�}���Y����[�^�D��e�d�d�e�f�l�G��I����V��B��U���d�l�u�k�u�m�F��I����V��^�D��e�d�d�d�u�}�W���H����X�^�D��d�d�e�d�f�m�G��H����V��NךU���g�`�h�u�g�l�F��H����W��_�E��d�d�d�d�{�W�W���K���F�_�D��d�d�d�e�g�l�F��I����W�d��U��l�u�k�w�g�l�F��H����V��^�D��d�e�e�w�w�}�W��@���D��_�D��d�e�e�e�f�m�F��H����D�=N��U��l�h�u�e�f�l�F��H����W��^�D��e�e�e�y�]�}�W��I���V��_�E��d�d�e�d�g�l�F��H����J�N��D��u�k�w�e�f�l�G��H����W��^�D��e�e�w�u�w�}�F��Y���V��_�D��e�e�e�d�g�l�F��H����FǻN��F��h�u�e�d�f�l�F��I����V��^�E��d�d�y�_�w�}�D��D���W��_�D��d�d�e�e�g�m�G��H���l�N�E���k�w�e�d�f�m�F��H����V��^�E��e�w�u�u�w�l�G���G����W��^�D��e�d�e�d�g�m�F��I���9F�_�B��u�e�d�d�f�l�F��H����V��^�D��d�y�_�u�w�n�O��Y����W��_�D��e�e�d�e�g�m�F��H���F�]�U��w�e�d�d�g�l�F��I����W��^�E��w�u�u�u�f�l�W���[����W��_�E��d�e�d�e�f�l�G��[��ƹF�_�H���e�d�d�d�f�l�G��H����V��^�E��y�_�u�u�d�o�J���I����W��_�D��d�e�e�e�f�m�G��U���F��]��K���e�d�d�e�f�l�F��I����V��_�D���u�u�u�d�f�}�I���I����V��_�D��d�d�e�d�g�l�G���Y���W��N��U��d�d�d�d�f�m�F��H����W��_�E���_�u�u�f�a�`�W��H����W��^�D��d�e�e�d�f�l�G��s���U��S�W��d�d�e�d�f�l�F��H����W��^�W���u�u�d�d�w�c�U��H����W��_�D��d�e�d�e�g�l�U���Y��� W��
P��E��d�d�d�d�f�m�G��I����V��^�Y�ߊu�u�f�e�j�}�G��H����W��^�D��e�e�d�e�g�m�[�ԜY����W�	N��E��d�e�d�d�g�m�F��H����W��_��U���u�d�g�u�i��G��H����W��^�E��e�d�d�e�g��W���Y���� F�L�D��d�d�d�d�g�l�G��I����V��L����u�f�a�h�w�m�F��H����W��_�D��e�e�e�d�g�q�}���Y����[�^�D��e�d�d�e�f�m�F��I����V��B��U���d�g�u�k�u�m�F��I����V��_�D��e�d�e�d�u�}�W���H����X�^�D��d�d�d�e�g�l�G��I����V��NךU���f�m�h�u�g�l�F��H����V��_�E��e�e�d�d�{�W�W���J���F�_�D��d�d�e�d�f�m�F��I����V�d��U��f�u�k�w�g�l�F��H����W��_�D��d�d�d�w�w�}�W��J���D��_�D��d�d�d�e�f�m�F��I����D�=N��U��g�h�u�e�f�l�F��H����V��_�D��e�d�d�y�]�}�W��J���V��_�E��d�e�e�d�f�m�F��H����J�N��D��u�k�w�e�f�l�G��H����V��_�E��e�d�w�u�w�}�F��Y���V��_�D��d�d�d�e�g�l�G��I����FǻN��F��h�u�e�d�f�l�F��H����W��_�D��d�d�y�_�w�}�D��D���W��_�D��e�d�e�e�g�m�F��H���l�N�F���k�w�e�d�f�m�F��I����W��^�E��d�w�u�u�w�l�D���G����W��^�D��d�d�e�e�f�m�G��H���9F�_�E��u�e�d�d�f�l�F��H����W��^�E��e�y�_�u�w�n�F��Y����W��_�D��d�d�d�e�f�l�G��H���F�]�U��w�e�d�d�g�l�F��I����W��^�D��w�u�u�u�f�i�W���[����W��_�D��e�d�e�e�g�l�F��[��ƹF�Z�H���e�d�d�d�f�l�F��I����V��_�D��y�_�u�u�d�h�J���I����W��_�D��e�e�e�e�f�m�G��U���F��X��K���e�d�d�e�f�l�F��I����V��_�D���u�u�u�d�c�}�I���I����V��_�E��d�e�e�e�g�m�G���Y���W��N��U��d�d�d�d�f�l�G��I����V��^�E���_�u�u�f�n�`�W��H����W��_�D��d�d�d�e�f�l�G��s���U��S�W��d�d�e�d�f�l�F��I����W��_�W���u�u�d�`�w�c�U��H����W��_�D��d�d�e�e�g�m�U���Y��� S��
P��E��d�d�d�d�f�m�F��H����W��_�Y�ߊu�u�f�f�j�}�G��H����W��^�D��d�e�d�e�g�m�[�ԜY����R�	N��E��d�e�d�d�f�m�G��I����V��_��U���u�d�`�u�i��G��H����W��^�D��e�d�d�d�f��W���Y����F�L�D��d�d�d�d�f�m�F��I����W��L����u�f�b�h�w�m�F��H����W��_�D��e�d�e�e�g�q�}���Y����[�^�D��e�d�d�d�g�l�G��I����V��B��U���d�`�u�k�u�m�F��I����W��_�D��e�e�d�e�u�}�W���H����X�^�D��d�d�d�d�g�m�G��H����W��NךU���f�d�h�u�g�l�F��H����W��^�E��d�e�d�e�{�W�W���J���F�_�D��d�d�d�d�f�m�F��H����V�d��U��c�u�k�w�g�l�F��H����W��_�D��d�e�d�w�w�}�W��O���D��_�D��d�d�d�d�g�m�G��H����D�=N��U��`�h�u�e�f�l�F��H����W��^�D��d�d�d�y�]�}�W��O���V��_�D��e�e�e�e�g�l�G��I����J�N��D��u�k�w�e�f�l�F��I����V��_�E��e�e�w�u�w�}�F��Y���V��_�E��e�e�e�d�f�l�G��I����FǻN��F��h�u�e�d�f�l�G��I����V��_�D��d�e�y�_�w�}�D��D���W��_�E��e�e�d�e�f�l�G��H���l�N�B���k�w�e�d�f�l�G��I����W��_�E��d�w�u�u�w�l�@���G����W��_�E��e�d�e�e�g�l�F��H���9F�_�F��u�e�d�d�f�m�G��I����V��_�D��e�y�_�u�w�n�C��Y����W��^�E��e�e�d�d�g�l�F��I���F�]�U��w�e�d�d�f�m�G��I����V��^�D��w�u�u�u�f�j�W���[����W��^�E��d�d�e�d�f�l�G��[��ƹF�Y�H���e�d�d�d�g�m�G��H����V��^�E��y�_�u�u�d�e�J���I����W��^�E��e�d�e�d�f�m�F��U���F�� W��K���e�d�d�d�g�m�G��I����W��^�D���u�u�u�d�o�}�I���I����W��^�E��d�d�d�d�f�m�G���Y���W��N��U��d�d�d�e�g�m�G��I����V��^�D���_�u�u�f�e�`�W��H����V��^�D��e�e�e�e�f�l�F��s���U��S�W��d�d�d�e�g�m�F��H����W��_�W���u�u�d�m�w�c�U��H����V��^�D��e�e�e�d�g�l�U���Y��� ^��
P��E��d�d�e�e�g�m�F��H����V��_�Y�ߊu�u�f�c�j�}�G��H����V��^�D��e�e�d�e�g�m�[�ԜY����Q�	N��E��d�d�e�e�g�l�F��H����W��^��U���u�d�m�u�i��G��H����V��_�D��e�e�e�d�g��W���Y����
F�L�D��d�e�e�e�f�m�G��I����V��L����u�f�e�h�w�m�F��H����V��^�D��d�d�e�e�f�q�}���Y����[�^�D��d�e�e�e�g�m�G��H����W��B��U���d�l�u�k�u�m�F��H����V��_�E��d�d�e�e�u�}�W���H����X�^�D��e�e�e�d�g�m�F��I����W��NךU���f�a�h�u�g�l�F��I����W��_�D��d�d�d�e�{�W�W���J���F�_�D��e�e�e�e�g�m�G��I����V�d��U��l�u�k�w�g�l�F��I����V��_�E��d�e�d�w�w�}�W��@���D��_�D��e�e�d�d�f�l�F��I����D�=N��U��m�h�u�e�f�l�F��I����W��^�E��e�e�d�y�]�}�W��@���V��_�D��e�e�e�d�f�m�G��I����J�N��D��u�k�w�e�f�l�F��I����W��_�D��d�d�w�u�w�}�F��Y���V��_�E��e�d�e�e�g�m�G��I����FǻN��A��h�u�e�d�f�l�G��I����V��_�D��d�e�y�_�w�}�C��D���W��_�E��e�d�e�d�g�m�F��H���l�N�E���k�w�e�d�f�l�G��I����V��_�D��e�w�u�u�w�l�G���G����W��_�E��d�e�e�d�f�l�G��H���9F�_�C��u�e�d�d�f�m�G��H����V��^�D��d�y�_�u�w�i�@��Y����W��^�E��d�e�e�d�g�m�G��I���F�Z�U��w�e�d�d�f�m�G��H����W��^�D��w�u�u�u�f�m�W���[����W��^�E��d�d�e�e�f�m�F��[��ƹF�_�H���e�d�d�d�g�m�G��H����W��^�D��y�_�u�u�c�l�J���I����W��^�E��d�d�d�e�f�m�G��U���F��\��K���e�d�d�d�g�m�G��H����V��^�E���u�u�u�d�f�}�I���I����W��^�E��e�e�d�d�f�m�F���Y���W��N��U��d�d�d�e�g�m�G��I����V��_�E���_�u�u�a�b�`�W��H����V��^�E��d�e�d�e�g�l�G��s���R��S�W��d�d�d�e�g�l�G��I����V��^�W���u�u�d�d�w�c�U��H����V��_�E��d�d�e�e�f�m�U���Y���W��
P��E��d�d�e�e�g�m�G��I����V��_�Y�ߊu�u�a�l�j�}�G��H����V��^�E��e�d�e�d�g�l�[�ԜY����V�	N��E��d�d�e�e�f�m�G��H����W��_��U���u�d�g�u�i��G��H����V��^�D��e�e�e�d�f��W���Y����F�L�D��d�e�e�e�g�l�G��I����W��L����u�a�f�h�w�m�F��H����V��_�D��d�e�e�e�f�q�}���Y����[�^�D��d�e�e�d�g�l�F��I����W��B��U���d�g�u�k�u�m�F��H����W��^�D��d�d�d�e�u�}�W���H����X�^�D��e�e�e�e�g�m�F��I����V��NךU���a�b�h�u�g�l�F��I����V��_�D��d�e�d�e�{�W�W���M���F�_�D��e�e�d�d�f�m�G��H����V�d��U��g�u�k�w�g�l�F��I����W��_�D��e�e�d�w�w�}�W��J���D��_�D��e�e�e�e�f�m�G��I����D�=N��U��d�h�u�e�f�l�F��I����W��_�E��d�d�e�y�]�}�W��K���V��_�D��e�d�d�e�g�m�G��I����J�N��D��u�k�w�e�f�l�F��I����V��_�D��d�e�w�u�w�}�F��Y���V��_�E��e�e�d�e�f�l�G��H����FǻN��A���h�u�e�d�f�l�G��I����W��^�D��d�e�y�_�w�}�C��D���W��_�E��d�d�d�d�f�l�F��I���l�N�F���k�w�e�d�f�l�G��H����V��_�E��e�w�u�u�w�l�D���G����W��_�E��d�e�d�e�g�l�F��I���9F�_�L��u�e�d�d�f�m�G��H����V��^�D��e�y�_�u�w�i�G��Y����W��^�E��e�d�e�e�f�m�G��I���F�Z�U��w�e�d�d�f�m�G��I����V��_�E��w�u�u�u�f�i�W���[����W��^�E��e�d�e�d�g�m�F��[��ƹF�Z�H���e�d�d�d�g�m�G��H����W��_�D��y�_�u�u�c�i�J���I����W��^�D��e�e�e�d�g�m�F��U���F��[��K���e�d�d�d�g�m�F��I����V��^�D���u�u�u�d�c�}�I���I����W��^�D��e�d�d�d�g�l�G���Y���W�� N��U��d�d�d�e�g�m�F��H����V��_�E���_�u�u�a�o�`�W��H����V��^�E��d�d�e�e�g�l�G��s���R��S�W��d�d�d�e�g�l�F��I����W��^�W���u�u�d�`�w�c�U��H����V��_�E��e�e�e�d�f�l�U���Y���S��
P��E��d�d�e�e�g�l�G��I����V��_�Y�ߊu�u�a�g�j�}�G��H����V��_�D��e�d�d�e�g�m�[�ԜY����U�	N��E��d�d�e�e�f�l�F��I����W��^��U���u�d�`�u�i��G��H����V��_�D��d�d�e�e�f��W���Y����F�L�D��d�e�e�e�f�l�G��H����V��L����u�a�c�h�w�m�F��H����V��_�E��d�e�d�d�g�q�}���Y����[�^�D��d�e�e�d�f�m�F��I����W��B��U���d�`�u�k�u�m�F��H����W��_�D��d�e�e�e�u�}�W���H����X�^�D��e�e�e�d�f�l�G��I����W��NךU���a�e�h�u�g�l�F��I����W��_�D��d�e�d�d�{�W�W���M���F�_�D��e�e�e�e�g�m�G��I����W�d��U��c�u�k�w�g�l�F��I����V��^�E��e�e�d�w�w�}�W��O���D��_�D��e�d�e�e�f�m�F��I����D�=N��U��a�h�u�e�f�l�F��I����V��_�D��d�e�e�y�]�}�W��L���V��_�D��e�e�e�d�g�m�G��H����J�N��D��u�k�w�e�f�l�F��I����W��_�E��d�e�w�u�w�}�F��Y���V��_�E��d�e�d�e�f�l�G��H����FǻN��A��h�u�e�d�f�l�G��H����W��^�E��e�d�y�_�w�}�C��D���W��_�E��e�e�e�d�f�l�F��I���l�N�B���k�w�e�d�f�l�G��I����V��_�D��e�w�u�u�w�l�@���G����W��_�E��e�d�d�e�g�m�G��H���9F�_�G��u�e�d�d�f�m�G��I����V��_�D��d�y�_�u�w�i�D��Y����W��^�E��d�e�e�e�g�l�F��I���F�Z�U��w�e�d�d�f�m�G��H����V��^�E��w�u�u�u�f�j�W���[����W��^�D��e�d�e�e�g�m�F��[��ƹF�Y�H���e�d�d�d�g�m�F��I����W��_�D��y�_�u�u�c�j�J���I����W��^�E��d�d�d�d�g�l�F��U���F�� V��K���e�d�d�d�g�m�G��H����V��^�E���u�u�u�d�`�}�I���I����W��^�E��e�d�d�e�g�l�G���Y���W��N��U��d�d�d�e�g�l�G��I����V��_�E���_�u�u�a�f�`�W��H����V��_�D��d�d�e�d�f�l�F��s���R��S�W��d�d�d�e�g�m�F��I����V��_�W���u�u�d�m�w�c�U��H����V��^�D��d�d�d�e�f�m�U���Y���^��
P��E��d�d�e�e�f�m�F��I����V��^�Y�ߊu�u�a�`�j�}�G��H����V��_�E��e�d�e�d�f�m�[�ԜY����P�	N��E��d�d�e�e�g�m�G��H����W��^��U���u�d�m�u�i��G��H����V��^�D��d�d�e�e�f��W���Y����F�L�D��d�e�e�d�f�m�G��I����W��L����u�a�l�h�w�m�F��H����W��^�D��d�d�d�e�f�q�}���Y����[�^�D��d�e�e�e�g�l�F��I����V��B��U���d�l�u�k�u�m�F��H����V��^�D��e�e�d�d�u�}�W���H����X�^�D��e�e�d�d�f�m�F��I����V��NךU���a�f�h�u�g�l�F��I����W��_�E��d�d�d�e�{�W�W���M���F�_�D��e�e�e�e�f�m�F��H����W�d��U��l�u�k�w�g�l�F��I����V��_�E��e�d�d�w�w�}�W��@���D��_�D��e�d�d�d�f�m�G��H����D�=N��U��b�h�u�e�f�l�F��I����V��^�E��d�e�e�y�]�}�W��A���V��_�D��e�e�d�e�f�m�F��I����J�N��D��u�k�w�e�f�l�F��I����V��^�E��e�e�w�u�w�}�F��Y���V��_�E��d�d�e�e�g�l�G��H����FǻN��@��h�u�e�d�f�l�G��H����V��_�E��e�e�y�_�w�}�B��D���W��_�E��e�d�d�d�g�m�F��H���l�N�E���k�w�e�d�f�l�G��I����V��_�E��e�w�u�u�w�l�G���G����W��_�E��d�d�e�d�f�m�F��H���9F�_�@��u�e�d�d�f�m�G��H����W��^�D��e�y�_�u�w�h�A��Y����W��^�E��d�d�e�d�g�m�G��H���F�[�U��w�e�d�d�f�m�G��H����V��^�D��w�u�u�u�f�m�W���[����W��^�D��d�d�d�d�f�l�G��[��ƹF�^�H���e�d�d�d�g�m�F��I����W��_�E��y�_�u�u�b�m�J���I����W��^�D��e�d�e�e�g�l�G��U���F��_��K���e�d�d�d�g�m�F��I����W��^�D���u�u�u�d�f�}�I���I����W��^�E��e�e�d�d�g�l�G���Y���W��N��U��d�d�d�e�g�l�G��I����W��_�D���_�u�u�`�c�`�W��H����V��_�E��e�d�e�d�f�m�F��s���S��S�W��d�d�d�e�g�l�G��I����W��_�W���u�u�d�d�w�c�U��H����V��_�D��e�d�d�e�g�l�U���Y���W��
P��E��d�d�e�e�f�m�F��H����V��^�Y�ߊu�u�`�m�j�}�G��H����V��^�D��e�e�d�d�f�l�[�ԜY����_�	N��E��d�d�e�e�f�m�F��H����W��^��U���u�d�g�u�i��G��H����V��^�D��d�d�e�e�g��W���Y����F�L�D��d�e�e�d�g�l�F��H����W��L����u�`�g�h�w�m�F��H����W��^�D��e�d�e�d�f�q�}���Y����[�^�D��d�e�e�d�f�m�G��H����W��B��U���d�g�u�k�u�m�F��H����W��^�D��d�d�e�d�u�}�W���H����X�^�D��e�e�d�e�g�m�G��H����V��NךU���`�c�h�u�g�l�F��I����V��_�E��e�d�d�d�{�W�W���L���F�_�D��e�e�d�d�f�l�F��I����W�d��U��g�u�k�w�g�l�F��I����W��_�D��e�e�e�w�w�}�W��K���D��_�D��e�d�e�d�f�m�F��H����D�=N��U���e�h�u�e�f�l�F��I����W��_�E��d�d�d�y�]�}�W��H���V��_�D��e�d�d�d�f�m�F��I����J�N��D��u�k�w�e�f�l�F��I����W��_�E��d�e�w�u�w�}�F��Y���V��_�E��d�e�d�d�f�l�G��I����FǻN��@��h�u�e�d�f�l�G��H����V��^�E��d�e�y�_�w�}�B��D���W��_�E��d�e�e�e�f�m�F��I���l�N�F���k�w�e�d�f�l�G��H����W��_�E��d�w�u�u�w�l�D���G����W��_�E��d�e�e�d�f�l�F��H���9F�_�M��u�e�d�d�f�m�G��H����V��_�E��e�y�_�u�w�h�N��Y����W��^�E��e�d�d�e�g�m�G��H���F�[�U��w�e�d�d�f�m�G��I����W��_�E��w�u�u�u�f�i�W���[����W��^�D��d�d�e�d�g�m�G��[��ƹF�Z�H���e�d�d�d�g�m�F��H����W��_�E��y�_�u�u�b�n�J���I����W��^�D��d�e�d�e�g�m�G��U���F��Z��K���e�d�d�d�g�m�F��H����V��_�D���u�u�u�d�c�}�I���I����W��^�D��d�e�e�d�f�m�G���Y���W��N��U��d�d�d�e�g�l�F��I����W��_�E���_�u�u�`�`�`�W��H����V��_�D��d�d�d�d�g�l�F��s���S��S�W��d�d�d�e�g�l�F��H����V��^�W���u�u�d�a�w�c�U��H����V��_�E��d�e�e�e�f�l�U���Y���S��
P��E��d�d�e�e�f�l�G��H����W��_�Y�ߊu�u�`�d�j�}�G��H����V��_�D��e�e�e�d�f�m�[�ԜY����T�	N��E��d�d�e�e�f�l�G��H����V��^��U���u�d�`�u�i��G��H����V��_�E��e�e�e�e�f��W���Y����F�L�D��d�e�e�d�f�l�F��I����V��L����u�`�`�h�w�m�F��H����W��_�E��d�d�e�d�f�q�}���Y����[�^�D��d�e�e�d�f�l�F��I����V��B��U���d�`�u�k�u�m�F��H����W��_�D��d�e�e�e�u�}�W���H����X�^�D��e�e�e�e�g�m�G��I����V��NךU���`�l�h�u�g�l�F��I����V��^�E��e�d�e�e�{�W�W���L���F�_�D��e�d�e�e�g�m�F��H����W�d��U��c�u�k�w�g�l�F��I����V��^�D��e�d�e�w�w�}�W��O���D��_�D��e�e�e�e�g�m�F��I����D�=N��U���f�h�u�e�f�l�F��I����V��_�E��d�d�e�y�]�}�W��M���V��_�D��d�e�e�e�g�m�G��H����J�N��D��u�k�w�e�f�l�F��H����V��_�D��d�d�w�u�w�}�F��Y���V��_�E��e�e�d�d�f�l�G��I����FǻN��@��h�u�e�d�f�l�G��I����W��_�E��e�d�y�_�w�}�B��D���W��_�E��e�e�d�d�g�l�F��H���l�N�C���k�w�e�d�f�l�G��I����V��^�E��e�w�u�u�w�l�@���G����W��_�E��e�d�d�d�g�m�F��I���9F�_�D��u�e�d�d�f�m�G��I����V��_�D��d�y�_�u�w�h�E��Y����W��^�D��d�e�e�d�g�m�G��H���F�[�U��w�e�d�d�f�m�F��H����V��_�D��w�u�u�u�f�j�W���[����W��^�E��e�e�e�e�g�m�F��[��ƹF�Y�H���e�d�d�d�g�m�G��I����V��_�D��y�_�u�u�b�k�J���I����W��^�E��d�d�e�d�f�m�G��U���F�� Y��K���e�d�d�d�g�l�G��I����V��_�E���u�u�u�d�`�}�I���I����W��_�E��d�e�d�d�g�m�G���Y���W��N��U��d�d�d�e�g�m�G��H����V��_�D���_�u�u�`�g�`�W��H����V��^�D��e�d�e�e�f�m�F��s���S��S�W��d�d�d�e�f�m�F��I����W��^�W���u�u�d�m�w�c�U��H����V��^�D��e�e�e�d�g�l�U���Y���^��
P��E��d�d�e�e�g�l�G��H����V��^�Y�ߊu�u�`�a�j�}�G��H����V��_�E��d�e�e�d�g�m�[�ԜY����S�	N��E��d�d�e�d�g�m�G��I����W��^��U���u�d�m�u�i��G��H����W��^�E��d�d�d�e�f��W���Y����F�L�D��d�e�e�e�f�m�G��I����V��L����u�`�m�h�w�m�F��H����V��^�D��d�e�d�e�g�q�}���Y����[�^�D��d�e�d�e�g�m�G��H����W��B��U���d�l�u�k�u�m�F��H����V��^�D��e�d�d�e�u�}�W���H����X�^�D��e�e�e�d�f�l�F��I����W��NךU���`�g�h�u�g�l�F��I����W��^�E��e�d�e�e�{�W�W���L���F�_�D��e�d�e�e�f�l�G��I����W�d��U��l�u�k�w�g�l�F��I����V��^�E��e�e�d�w�w�}�W��@���D��_�D��e�e�d�e�g�m�G��I����D�=N��U���c�h�u�e�f�l�F��I����V��^�D��e�d�e�y�]�}�W��N���V��_�D��d�e�d�e�g�m�G��H����J�N��D��u�k�w�e�f�l�F��H����V��_�E��d�d�w�u�w�}�F��Y���V��_�E��e�d�e�e�g�l�F��H����FǻN��C��h�u�e�d�f�l�G��I����W��^�E��e�e�y�_�w�}�A��D���W��_�E��e�d�d�d�f�m�G��H���l�N�E���k�w�e�d�f�l�G��I����W��_�E��e�w�u�u�w�l�G���G����W��_�E��d�d�d�e�g�l�G��I���9F�_�A��u�e�d�d�f�m�G��H����W��^�D��e�y�_�u�w�k�B��Y����W��^�D��d�d�e�d�g�l�F��I���F�X�U��w�e�d�d�f�m�F��H����V��_�D��w�u�u�u�f�m�W���[����W��^�E��d�d�e�d�f�m�F��[��ƹF�^�H���e�d�d�d�g�m�G��I����V��^�D��y�_�u�u�a�d�J���I����W��^�D��e�e�e�e�f�m�G��U���F��^��K���e�d�d�d�g�l�F��I����W��_�D���u�u�u�d�f�}�I���I����W��_�E��e�d�e�d�g�l�G���Y���W��N��U��d�d�d�e�g�m�G��I����V��_�E���_�u�u�c�d�`�W��H����V��^�E��d�e�e�d�f�m�G��s���P��S�W��d�d�d�e�f�l�G��I����W��^�W���u�u�d�d�w�c�U��H����V��_�D��d�d�d�e�g�l�U���Y���W��
P��E��d�d�e�e�g�m�F��I����W��^�Y�ߊu�u�c�b�j�}�G��H����V��^�D��d�e�e�e�f�m�[�ԜY����^�	N��E��d�d�e�d�f�m�F��I����V��_��U���u�d�d�u�i��G��H����W��^�D��e�d�e�e�f��W���Y����F�L�D��d�e�e�e�g�m�G��H����V��L����u�c�d�h�w�m�F��H����V��^�D��e�d�d�e�f�q�}���Y����[�^�D��d�e�d�d�f�m�G��I����V��B��U���d�g�u�k�u�m�F��H����W��^�D��e�e�d�e�u�}�W���H����X�^�D��e�e�e�e�g�m�G��H����W��NךU���c�`�h�u�g�l�F��I����V��_�E��e�e�e�d�{�W�W���O���F�_�D��e�d�d�d�f�l�F��I����V�d��U��g�u�k�w�g�l�F��I����W��_�E��d�d�d�w�w�}�W��K���D��_�D��e�e�e�d�f�m�G��I����D�=N��U��l�h�u�e�f�l�F��I����W��_�D��d�d�d�y�]�}�W��I���V��_�D��d�d�d�d�g�l�G��H����J�N��D��u�k�w�e�f�l�F��H����W��^�E��d�d�w�u�w�}�F��Y���V��_�E��e�e�d�d�g�l�F��H����FǻN��C��h�u�e�d�f�l�G��I����V��_�E��d�d�y�_�w�}�A��D���W��_�E��d�e�e�d�f�l�G��I���l�N�F���k�w�e�d�f�l�G��H����W��_�D��d�w�u�u�w�l�D���G����W��_�E��d�e�e�d�g�m�G��H���9F�_�B��u�e�d�d�f�m�G��H����W��_�D��d�y�_�u�w�k�O��Y����W��^�D��e�d�d�e�g�l�F��I���F�X�U��w�e�d�d�f�m�F��I����W��_�D��w�u�u�u�f�i�W���[����W��^�E��d�e�d�e�f�m�F��[��ƹF�Z�H���e�d�d�d�g�m�G��H����V��_�E��y�_�u�u�a�o�J���I����W��^�D��d�e�e�e�f�m�G��U���F��]��K���e�d�d�d�g�l�F��H����V��_�E���u�u�u�d�c�}�I���I����W��_�D��d�d�d�d�g�l�F���Y���W��N��U��d�d�d�e�g�m�F��H����V��_�D���_�u�u�c�a�`�W��H����V��^�D��d�e�d�d�f�l�G��s���P��S�W��d�d�d�e�f�l�F��I����V��_�W���u�u�d�a�w�c�U��H����V��_�E��d�e�e�e�g�l�U���Y���R��
P��E��d�d�e�e�g�l�G��I����V��_�Y�ߊu�u�c�e�j�}�G��H����V��_�D��d�e�e�d�g�l�[�ԜY����W�	N��E��d�d�e�d�f�l�F��I����W��^��U���u�d�`�u�i��G��H����W��_�E��e�e�e�d�g��W���Y���� F�L�D��d�e�e�e�f�l�F��I����W��L����u�c�a�h�w�m�F��H����V��_�D��d�e�d�e�g�q�}���Y����[�^�D��d�e�d�d�f�l�G��H����W��B��U���d�`�u�k�u�m�F��H����W��_�D��e�e�e�d�u�}�W���H����X�^�D��e�e�e�d�f�l�G��I����V��NךU���c�m�h�u�g�l�F��I����V��^�D��e�e�d�d�{�W�W���O���F�_�D��e�d�e�e�g�l�G��I����V�d��U��c�u�k�w�g�l�F��I����V��^�D��d�e�e�w�w�}�W��O���D��_�D��e�d�e�e�g�m�F��H����D�=N��U��g�h�u�e�f�l�F��I����V��^�D��d�d�d�y�]�}�W��J���V��_�D��d�e�e�d�g�m�F��I����J�N��D��u�k�w�e�f�l�F��H����W��_�D��e�e�w�u�w�}�F��Y���V��_�E��d�e�d�e�g�l�F��H����FǻN��C��h�u�e�d�f�l�G��H����W��^�E��d�d�y�_�w�}�A��D���W��_�E��e�e�e�d�f�m�F��I���l�N�C���k�w�e�d�f�l�G��I����W��^�D��d�w�u�u�w�l�A���G����W��_�E��e�d�d�e�g�l�G��I���9F�_�E��u�e�d�d�f�m�G��I����W��_�E��e�y�_�u�w�k�F��Y����W��^�D��d�e�e�d�g�l�G��H���F�X�U��w�e�d�d�f�m�F��H����V��^�D��w�u�u�u�f�j�W���[����W��^�D��e�d�e�e�g�l�G��[��ƹF�Y�H���e�d�d�d�g�m�F��I����V��^�D��y�_�u�u�a�h�J���I����W��^�E��d�d�d�d�f�l�F��U���F�� X��K���e�d�d�d�g�l�G��H����W��_�E���u�u�u�d�`�}�I���I����W��_�E��e�e�e�d�f�m�G���Y���W��N��U��d�d�d�e�g�l�G��I����W��_�D���_�u�u�c�n�`�W��H����V��_�D��e�d�d�d�g�l�F��s���P��S�W��d�d�d�e�f�m�F��I����V��^�W���u�u�d�m�w�c�U��H����V��^�D��e�d�e�e�f�m�U���Y���^��
P��E��d�d�e�e�f�m�F��H����W��_�Y�ߊu�u�c�f�j�}�G��H����V��^�D��d�e�d�e�g�m�[�ԜY����R�	N��E��d�d�e�d�g�m�G��I����W��_��U���u�d�m�u�i��G��H����W��^�D��d�e�d�e�f��W���Y����F�L�D��d�e�e�d�f�m�F��H����V��L����u�c�b�h�w�m�F��H����W��^�E��e�e�e�d�g�q�}���Y����[�^�D��d�e�d�e�g�l�G��I����V��B��U���d�m�u�k�u�m�F��H����V��_�E��d�e�d�d�u�}�W���H����X�^�D��e�e�d�d�f�m�F��H����V��NךU���c�d�h�u�g�l�F��I����W��^�D��e�d�e�d�{�W�W���O���F�_�D��e�d�e�e�g�l�G��I����V�d��U��l�u�k�w�g�l�F��I����V��^�D��d�d�d�w�w�}�W��@���D��_�D��e�d�d�d�g�l�F��I����D�=N��U��`�h�u�e�f�l�F��I����W��_�E��e�d�e�y�]�}�W��O���V��_�D��d�e�d�e�g�m�G��I����J�N��D��u�k�w�e�f�l�F��H����V��_�D��e�e�w�u�w�}�F��Y���V��_�E��d�d�e�d�f�l�F��I����FǻN��C��h�u�e�d�f�l�G��H����W��_�D��e�e�y�_�w�}�@��D���W��_�E��e�d�d�d�g�m�G��I���l�N�E���k�w�e�d�f�l�G��I����V��^�D��e�w�u�u�w�l�G���G����W��_�E��d�e�d�d�f�l�F��I���9F�_�F��u�e�d�d�f�m�G��H����W��_�E��e�y�_�u�w�j�C��Y����W��^�D��d�e�e�e�g�m�F��H���F�Y�U��w�e�d�d�f�m�F��H����W��^�D��w�u�u�u�f�m�W���[����W��^�D��d�e�d�d�g�l�F��[��ƹF� ^�H���e�d�d�d�g�m�F��H����W��_�D��y�_�u�u�`�e�J���I����W��^�E��d�d�e�e�f�l�F��U���F��W��K���e�d�d�d�g�l�F��I����V��^�E���u�u�u�d�f�}�I���I����W��_�E��e�d�d�e�f�l�G���Y���W��N��U��d�d�d�e�g�l�G��H����V��^�D���_�u�u�b�e�`�W��H����V��_�E��e�e�e�e�g�l�G��s���Q��S�W��d�d�d�e�f�l�G��H����W��_�W���u�u�d�d�w�c�U��H����V��_�E��d�e�d�e�f�l�U���Y���W��
P��E��d�d�e�e�f�m�G��H����W��_�Y�ߊu�u�b�c�j�}�G��H����V��^�E��e�d�e�e�g�m�[�ԜY����Q�	N��E��d�d�e�d�f�m�G��H����V��_��U���u�d�d�u�i��G��H����W��^�D��e�e�d�e�f��W���Y����
F�L�D��d�e�e�d�g�l�G��I����V��L����u�b�e�h�w�m�F��H����W��_�E��d�e�d�d�f�q�}���Y����[�^�D��d�e�d�d�g�l�F��I����V��B��U���d�g�u�k�u�m�F��H����W��^�D��d�e�e�e�u�}�W���H����X�^�D��e�e�d�e�g�m�F��H����V��NךU���b�a�h�u�g�l�F��I����V��_�E��e�e�d�e�{�W�W���N���F�_�D��e�d�d�d�f�m�F��H����V�d��U��g�u�k�w�g�l�F��I����W��_�E��d�d�d�w�w�}�W��K���D��_�D��e�d�e�e�f�l�G��I����D�=N��U��m�h�u�e�f�l�F��I����V��_�D��d�e�d�y�]�}�W��@���V��_�D��d�d�d�e�f�m�F��I����J�N��D��u�k�w�e�f�l�F��H����V��_�E��d�d�w�u�w�}�F��Y���V��_�E��d�e�d�d�f�l�G��H����FǻN��B��h�u�e�d�f�l�G��H����V��_�E��d�e�y�_�w�}�@��D���W��_�E��d�d�d�e�g�m�F��H���l�N�F���k�w�e�d�f�l�G��H����W��^�E��d�w�u�u�w�l�D���G����W��_�E��d�e�e�d�f�m�G��I���9F�_�C��u�e�d�d�f�m�G��H����W��^�E��e�y�_�u�w�j�@��Y����W��^�D��e�e�d�e�f�l�G��I���F�Y�U��w�e�d�d�f�m�F��I����W��^�E��w�u�u�u�f�n�W���[����W��^�D��e�e�d�e�g�l�F��[��ƹF� Z�H���e�d�d�d�g�m�F��I����V��_�D��y�_�u�u�`�l�J���I����W��^�D��e�e�e�e�f�m�G��U���F��\��K���e�d�d�d�g�l�F��I����V��_�D���u�u�u�d�c�}�I���I����W��_�D��d�d�e�e�g�l�G���Y���W��N��U��d�d�d�e�g�l�F��H����V��^�E���_�u�u�b�b�`�W��H����V��_�E��e�d�d�d�g�m�F��s���Q��S�W��d�d�d�e�f�l�G��I����W��_�W���u�u�d�a�w�c�U��H����V��_�D��e�d�e�d�g�l�U���Y���R��
P��E��d�d�e�e�f�l�G��H����W��^�Y�ߊu�u�b�l�j�}�G��H����V��_�E��d�e�e�d�f�m�[�ԜY����V�	N��E��d�d�e�d�f�l�G��I����V��_��U���u�d�`�u�i��G��H����W��_�E��e�d�d�e�f��W���Y����F�L�D��d�e�e�d�f�m�G��I����W��L����u�b�f�h�w�m�F��H����W��^�E��d�d�e�e�g�q�}���Y����[�^�D��d�e�d�d�f�m�G��I����V��B��U���d�`�u�k�u�m�F��H����W��^�E��d�e�d�d�u�}�W���H����X�^�D��e�e�d�d�f�l�F��I����V��NךU���b�b�h�u�g�l�F��I����W��_�E��d�e�d�e�{�W�W���N���F�_�D��e�d�d�d�f�m�F��I����W�d��U��`�u�k�w�g�l�F��I����W��^�D��d�d�d�w�w�}�W��O���D��_�D��e�d�d�d�f�m�F��I����D�=N��U��d�h�u�e�f�l�F��H����V��_�E��e�e�d�y�]�}�W��K���V��_�D��e�e�e�e�f�l�G��I����J�N��D��u�k�w�e�f�l�F��I����V��^�D��e�e�w�u�w�}�F��Y���V��_�E��e�e�e�e�g�m�G��H����FǻN��B���h�u�e�d�f�l�G��I����V��^�D��d�e�y�_�w�}�@��D���W��_�E��e�e�d�e�f�m�F��I���l�N�C���k�w�e�d�f�l�G��I����V��^�E��e�w�u�u�w�l�A���G����W��_�D��e�d�e�e�f�l�G��H���9F�_�L��u�e�d�d�f�m�F��I����V��^�E��d�y�_�u�w�j�G��Y����W��^�E��e�e�d�e�g�m�F��I���F�Y�U��w�e�d�d�f�m�G��I����W��_�E��w�u�u�u�f�j�W���[����W��^�E��d�d�e�e�f�m�G��[��ƹF� Y�H���e�d�d�d�g�l�G��H����V��^�D��y�_�u�u�`�i�J���I����W��_�E��e�e�e�e�f�m�G��U���F�� [��K���e�d�d�d�g�m�G��I����V��_�E���u�u�u�d�`�}�I���I����W��^�E��d�d�d�d�f�l�G���Y���W�� N��U��d�d�d�e�f�m�G��I����V��_�E���_�u�u�b�o�`�W��H����V��^�D��d�d�d�e�g�m�F��s���Q��S�W��d�d�d�e�g�m�F��I����V��_�W���u�u�d�m�w�c�U��H����V��^�E��d�d�e�e�g�l�U���Y���^��
P��E��d�d�e�d�g�m�F��I����V��_�Y�ߊu�u�b�g�j�}�G��H����W��^�E��d�d�e�e�f�m�[�ԜY����U�	N��E��d�d�e�e�g�l�G��I����V��^��U���u�d�m�u�i��G��H����V��_�E��d�d�d�d�f��W���Y����F�L�D��d�e�d�e�g�l�G��H����V��L����u�b�c�h�w�m�F��H����V��_�D��e�d�e�d�g�q�}���Y����[�^�D��d�e�e�e�g�m�G��I����V��B��U���d�m�u�k�u�m�F��H����V��^�D��d�e�e�d�u�}�W���H����X�^�D��e�d�e�d�g�l�F��I����W��NךU���b�e�h�u�g�l�F��I����W��^�E��e�d�e�d�{�W�W���N���F�_�D��e�e�e�e�f�l�F��I����W�d��U��l�u�k�w�g�l�F��I����V��^�D��e�d�e�w�w�}�W��@���D��_�D��d�e�d�e�f�l�F��I����D�=N��U��a�h�u�e�f�l�F��H����W��_�E��d�e�d�y�]�}�W��L���V��_�D��e�e�e�e�g�m�F��H����J�N��D��u�k�w�e�f�l�F��I����V��_�E��e�d�w�u�w�}�F��Y���V��_�E��e�d�d�e�f�m�F��H����FǻN��B��h�u�e�d�f�l�G��I����V��^�E��d�e�y�_�w�}�@��D���W��_�E��e�e�d�e�f�l�F��I���l�N�E���k�w�e�d�f�l�G��I����V��^�E��d�w�u�u�w�l�G���G����W��_�D��d�e�e�e�f�m�F��H���9F�_�G��u�e�d�d�f�m�F��H����W��_�D��e�y�_�u�w�e�D��Y����W��^�E��d�e�d�d�g�l�G��H���F�V�U��w�e�d�d�f�m�G��H����V��_�D��w�u�u�u�f�m�W���[����W��^�E��e�d�e�d�f�l�G��[��ƹF�^�H���e�d�d�d�g�l�G��I����W��_�D��y�_�u�u�o�j�J���I����W��_�E��e�e�e�e�f�l�F��U���F��V��K���e�d�d�d�g�m�G��I����W��^�E���u�u�u�d�g�}�I���I����W��^�D��d�e�e�d�f�l�G���Y���W��N��U��d�d�d�e�f�m�F��I����V��_�D���_�u�u�m�f�`�W��H����V��^�D��d�d�d�e�f�l�F��s���^��S�W��d�d�d�e�g�m�F��I����W��_�W���u�u�d�d�w�c�U��H����V��^�D��d�d�e�d�f�l�U���Y���W��
P��E��d�d�e�d�g�m�G��I����V��_�Y�ߊu�u�m�`�j�}�G��H����W��^�E��d�e�d�d�g�l�[�ԜY����P�	N��E��d�d�e�e�f�m�G��I����W��^��U���u�d�d�u�i��G��H����V��^�E��d�e�d�e�g��W���Y����F�L�D��d�e�d�e�g�m�G��H����V��L����u�m�l�h�w�m�F��H����V��^�D��d�d�e�e�g�q�}���Y����[�^�D��d�e�e�d�g�m�G��H����W��B��U���d�g�u�k�u�m�F��H����W��^�D��e�d�d�e�u�}�W���H����X�^�D��e�d�e�e�f�l�F��H����V��NךU���m�f�h�u�g�l�F��I����V��_�D��d�e�e�d�{�W�W���A���F�_�D��e�e�d�e�f�l�G��I����W�d��U��g�u�k�w�g�l�F��I����V��^�E��e�d�d�w�w�}�W��K���D��_�D��d�e�e�d�f�l�G��I����D�=N��U��b�h�u�e�f�l�F��H����V��_�D��e�d�d�y�]�}�W��A���V��_�D��e�d�d�e�f�l�F��I����J�N��D��u�k�w�e�f�l�F��I����V��^�E��d�e�w�u�w�}�F��Y���V��_�E��e�e�e�e�g�m�G��H����FǻN��M��h�u�e�d�f�l�G��I����V��^�E��e�d�y�_�w�}�O��D���W��_�E��d�d�d�e�g�l�F��I���l�N�F���k�w�e�d�f�l�G��H����W��^�D��e�w�u�u�w�l�D���G����W��_�D��e�d�e�e�f�m�F��I���9F�_�@��u�e�d�d�f�m�F��I����V��^�E��e�y�_�u�w�e�A��Y����W��^�E��d�e�d�e�g�l�F��H���F�V�U��w�e�d�d�f�m�G��H����V��^�D��w�u�u�u�f�n�W���[����W��^�E��d�e�d�d�f�m�G��[��ƹF�]�H���e�d�d�d�g�l�G��H����V��_�E��y�_�u�u�o�m�J���I����W��_�D��e�e�d�d�g�m�G��U���F��_��K���e�d�d�d�g�m�F��I����V��^�D���u�u�u�d�c�}�I���I����W��^�D��d�d�d�e�g�l�F���Y���W��N��U��d�d�d�e�f�m�F��H����V��_�E���_�u�u�m�c�`�W��H����V��^�E��d�e�d�e�g�l�G��s���^��S�W��d�d�d�e�g�l�G��I����V��_�W���u�u�d�a�w�c�U��H����V��_�E��e�d�d�d�g�l�U���Y���R��
P��E��d�d�e�d�g�l�F��H����V��_�Y�ߊu�u�m�m�j�}�G��H����W��_�E��d�d�d�e�g�l�[�ԜY����_�	N��E��d�d�e�e�f�m�G��I����W��_��U���u�d�`�u�i��G��H����V��^�E��e�e�e�d�f��W���Y����F�L�D��d�e�d�e�f�l�G��H����W��L����u�m�g�h�w�m�F��H����V��_�E��e�e�e�e�g�q�}���Y����[�^�D��d�e�e�d�g�l�F��H����W��B��U���d�`�u�k�u�m�F��H����W��^�E��e�e�e�d�u�}�W���H����X�^�D��e�d�e�d�g�l�G��I����V��NךU���m�c�h�u�g�l�F��I����W��_�D��d�d�d�e�{�W�W���A���F�_�D��e�e�d�d�f�m�G��H����W�d��U��`�u�k�w�g�l�F��I����W��_�E��d�e�d�w�w�}�W��L���D��_�D��d�e�d�e�f�l�F��H����D�=N��U��e�h�u�e�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H���V��_�D��e�d�d�e�f�l�F��I����J�N��D��u�k�w�e�f�l�F��I����V��^�E��d�e�w�u�w�}�F��Y���V��_�E��e�d�d�d�f�l�G��I����FǻN��M��h�u�e�d�f�l�G��I����V��_�D��e�d�y�_�w�}�O��D���W��_�E��d�d�d�e�g�l�F��I���l�N�C���k�w�e�d�f�l�G��H����W��^�E��e�w�u�u�w�l�A���G����W��_�D��e�e�e�e�f�m�G��H���9F�_�M��u�e�d�d�f�m�F��I����W��^�E��e�y�_�u�w�e�N��Y����W��^�E��e�e�e�d�f�m�F��I���F�V�U��w�e�d�d�f�m�G��I����V��^�E��w�u�u�u�f�j�W���[����W��^�D��e�e�e�d�g�m�G��[��ƹF�Y�H���e�d�d�d�g�l�F��I����W��^�D��y�_�u�u�o�n�J���I����W��_�E��d�d�e�e�f�l�G��U���F�� Z��K���e�d�d�d�g�m�G��I����W��_�D���u�u�u�d�`�}�I���I����W��^�E��e�d�d�d�g�l�G���Y���W��N��U��d�d�d�e�f�l�G��H����W��^�E���_�u�u�m�`�`�W��H����V��_�E��e�d�e�e�f�l�F��s���^��S�W��d�d�d�e�g�m�G��H����W��_�W���u�u�d�b�w�c�U��H����V��^�D��d�d�e�e�f�l�U���Y���^��
P��E��d�d�e�d�f�m�F��H����V��^�Y�ߊu�u�m�d�j�}�G��H����W��^�E��e�e�e�e�g�l�[�ԜY����T�	N��E��d�d�e�e�g�l�G��I����V��^��U���u�d�m�u�i��G��H����V��_�D��e�d�e�d�g��W���Y����F�L�D��d�e�d�d�g�m�G��I����W��L����u�m�`�h�w�m�F��H����W��^�D��d�e�d�e�f�q�}���Y����[�^�D��d�e�e�e�f�l�G��I����V��B��U���d�m�u�k�u�m�F��H����V��^�E��e�e�e�e�u�}�W���H����X�^�D��e�d�d�e�f�m�G��I����V��NךU���m�l�h�u�g�l�F��I����V��_�D��d�e�e�e�{�W�W���A���F�_�D��e�e�e�d�g�l�G��I����W�d��U��l�u�k�w�g�l�F��I����W��^�E��e�d�e�w�w�}�W��@���D��_�D��d�d�e�d�g�l�F��I����D�=N��U��f�h�u�e�f�l�F��H����W��^�E��e�d�e�y�]�}�W��M���V��_�D��e�e�e�e�g�l�G��I����J�N��D��u�k�w�e�f�l�F��I����V��_�D��d�e�w�u�w�}�F��Y���V��_�E��d�d�e�d�f�l�F��I����FǻN��M��h�u�e�d�f�l�G��H����W��^�D��d�e�y�_�w�}�O��D���W��_�E��e�e�d�d�g�m�G��I���l�N�L���k�w�e�d�f�l�G��I����V��^�E��e�w�u�u�w�l�G���G����W��_�D��d�e�d�e�g�l�G��H���9F�_�D��u�e�d�d�f�m�F��H����W��^�E��d�y�_�u�w�d�E��Y����W��^�E��e�e�d�e�f�m�G��H���F�W�U��w�e�d�d�f�m�G��I����W��_�E��w�u�u�u�f�m�W���[����W��^�D��d�e�e�e�f�m�G��[��ƹF�^�H���e�d�d�d�g�l�F��H����W��_�E��y�_�u�u�n�k�J���I����W��_�E��d�e�d�d�f�l�G��U���F��Y��K���e�d�d�d�g�m�G��H����V��^�D���u�u�u�d�g�}�I���I����W��^�D��e�d�d�e�g�l�F���Y���W��N��U��d�d�d�e�f�l�F��I����V��_�E���_�u�u�l�g�`�W��H����V��_�D��d�e�e�e�f�l�G��s���_��S�W��d�d�d�e�g�m�F��I����W��_�W���u�u�d�d�w�c�U��H����V��^�E��e�d�e�e�f�l�U���Y���
W��
P��E��d�d�e�d�f�l�G��H����V��_�Y�ߊu�u�l�a�j�}�G��H����W��_�D��e�d�d�d�g�m�[�ԜY����S�	N��E��d�d�e�e�g�l�G��H����W��_��U���u�d�d�u�i��G��H����V��_�D��e�d�d�d�f��W���Y����F�L�D��d�e�d�d�f�l�F��H����V��L����u�l�m�h�w�m�F��H����W��_�E��e�e�e�e�g�q�}���Y����[�^�D��d�e�e�e�f�l�F��I����V��B��U���d�g�u�k�u�m�F��H����V��_�D��e�e�d�d�u�}�W���H����X�^�D��e�d�d�d�f�l�F��H����V��NךU���l�g�h�u�g�l�F��I����V��^�E��e�e�d�d�{�W�W���@���F�_�D��e�e�d�e�g�m�G��I����V�d��U��g�u�k�w�g�l�F��I����V��_�E��d�d�e�w�w�}�W��K���D��_�D��d�d�e�e�g�l�G��I����D�=N��U��c�h�u�e�f�l�F��H����V��_�E��e�d�d�y�]�}�W��N���V��_�D��e�d�e�d�g�l�F��H����J�N��D��u�k�w�e�f�l�F��I����V��^�E��d�d�w�u�w�}�F��Y���V��_�E��d�e�d�e�g�l�F��I����FǻN��L��h�u�e�d�f�l�G��H����W��^�E��d�d�y�_�w�}�N��D���W��_�E��d�e�e�d�f�l�G��H���l�N�F���k�w�e�d�f�l�G��H����V��^�E��e�w�u�u�w�l�D���G����W��_�D��e�d�e�d�g�l�G��I���9F�_�A��u�e�d�d�f�m�F��I����W��^�D��d�y�_�u�w�d�B��Y����W��^�E��d�e�e�e�f�l�G��I���F�W�U��w�e�d�d�f�m�G��H����W��_�D��w�u�u�u�f�n�W���[����W��^�D��e�d�e�d�f�l�F��[��ƹF�]�H���e�d�d�d�g�l�F��I����V��_�D��y�_�u�u�n�d�J���I����W��_�D��d�e�e�d�f�l�G��U���F��^��K���e�d�d�d�g�m�F��H����V��^�D���u�u�u�d�c�}�I���I����W��^�E��d�e�e�d�f�l�G���Y���W��N��U��d�d�d�e�f�l�G��I����V��^�D���_�u�u�l�d�`�W��H����V��_�D��d�d�d�d�g�m�F��s���_��S�W��d�d�d�e�g�l�F��I����W��^�W���u�u�d�a�w�c�U��H����V��_�D��d�d�d�e�g�m�U���Y���
R��
P��E��d�d�e�d�f�m�F��H����V��^�Y�ߊu�u�l�b�j�}�G��H����W��^�D��d�d�e�d�g�m�[�ԜY����^�	N��E��d�d�e�e�f�l�F��I����V��_��U���u�d�a�u�i��G��H����V��^�E��e�d�e�d�g��W���Y����F�L�D��d�e�d�d�f�m�G��H����V��L����u�l�d�h�w�m�F��H����W��^�E��d�d�d�e�f�q�}���Y����[�^�D��d�e�e�d�g�m�F��H����W��B��U���d�`�u�k�u�m�F��H����W��_�D��e�e�e�d�u�}�W���H����X�^�D��e�d�d�d�g�l�G��H����W��NךU���l�`�h�u�g�l�F��I����W��_�E��e�d�d�e�{�W�W���@���F�_�D��e�e�d�e�g�m�F��H����V�d��U��`�u�k�w�g�l�F��I����V��_�D��e�d�d�w�w�}�W��L���D��_�D��d�d�d�d�f�l�F��H����D�=N��U��l�h�u�e�f�l�F��H����W��_�E��d�e�e�y�]�}�W��I���V��_�D��e�d�e�d�g�l�G��H����J�N��D��u�k�w�e�f�l�F��I����W��^�E��e�d�w�u�w�}�F��Y���V��_�E��d�d�d�d�g�l�F��H����FǻN��L��h�u�e�d�f�l�G��H����V��_�E��d�d�y�_�w�}�N��D���W��_�E��d�d�e�d�g�m�F��I���l�N�C���k�w�e�d�f�l�G��H����V��^�D��e�w�u�u�w�l�A���G����W��_�D��d�e�d�d�g�m�G��H���9F�_�B��u�e�d�d�f�m�F��H����W��^�D��d�y�_�u�w�d�O��Y����W��^�E��d�d�e�e�f�m�G��H���F�W�U��w�e�d�d�f�m�G��H����V��_�E��w�u�u�u�f�j�W���[����W��^�D��d�e�e�d�g�l�F��[��ƹF�Y�H���e�d�d�d�g�l�F��H����V��^�E��y�_�u�u�n�o�J���I����W��_�D��e�e�e�e�f�l�G��U���F�� ]��K���e�d�d�d�g�m�F��I����W��_�D���u�u�u�d�`�}�I���I����W��^�D��e�d�d�e�f�m�G���Y���W��N��U��d�d�d�e�f�l�F��H����W��^�E���_�u�u�l�a�`�W��H����V��_�D��d�e�d�d�g�l�G��s���_��S�W��d�d�d�e�f�m�G��I����V��_�W���u�u�d�b�w�c�U��H����V��^�E��d�e�e�d�g�m�U���Y���
Q��
P��E��d�d�e�d�g�m�G��H����W��_�Y�ߊu�u�l�e�j�}�G��H����W��^�E��d�e�d�d�f�m�[�ԜY����W�	N��E��d�d�e�d�g�m�F��H����W��^��U���u�d�m�u�i��G��H����W��^�D��e�e�e�e�g��W���Y���� F�L�D��d�e�d�e�g�m�F��H����V��L����u�l�a�h�w�m�F��H����V��_�E��d�e�d�e�f�q�}���Y����[�^�D��d�e�d�e�g�m�F��H����W��B��U���d�m�u�k�u�m�F��H����V��^�D��e�e�d�d�u�}�W���H����X�^�D��e�d�e�e�f�l�F��I����W��NךU���l�m�h�u�g�l�F��I����V��^�D��d�d�d�e�{�W�W���@���F�_�D��e�d�e�e�f�m�G��I����V�d��U��l�u�k�w�g�l�F��I����V��_�D��e�e�d�w�w�}�W��@���D��_�D��d�e�e�e�g�m�G��H����D�=N��U��g�h�u�e�f�l�F��H����V��^�D��e�e�e�y�]�}�W��J���V��_�D��d�e�d�e�g�m�F��I����J�N��D��u�k�w�e�f�l�F��H����V��^�E��d�d�w�u�w�}�F��Y���V��_�E��e�e�e�e�f�m�F��H����FǻN��L��h�u�e�d�f�l�G��I����V��_�E��d�d�y�_�w�}�N��D���W��_�E��e�d�d�d�g�l�F��H���l�N�L���k�w�e�d�f�l�G��I����V��_�D��e�w�u�u�w�l�N���G����W��_�D��e�d�e�e�f�m�G��I���9F�\�E��u�e�d�d�f�m�F��I����W��^�D��d�y�_�u�w�m�F��Y����W��^�D��d�e�d�e�g�m�F��H���F�^�U��w�e�d�d�f�m�F��H����W��_�D��w�u�u�u�e�m�W���[����W��^�E��d�e�d�d�g�m�F��[��ƹF�^�H���e�d�d�d�g�l�G��H����V��_�E��y�_�u�u�g�h�J���I����W��_�E��e�e�e�e�g�m�G��U���F��X��K���e�d�d�d�g�l�G��I����V��_�E���u�u�u�g�g�}�I���I����W��_�D��d�e�d�d�g�l�F���Y���T��N��U��d�d�d�e�f�m�F��H����W��_�E���_�u�u�e�n�`�W��H����V��^�E��e�e�e�e�f�l�G��s���V��S�W��d�d�d�e�f�m�G��H����V��_�W���u�u�g�d�w�c�U��H����V��^�E��d�d�d�e�g�l�U���Y���W��
P��E��d�d�e�d�g�l�F��I����V��_�Y�ߊu�u�e�f�j�}�G��H����W��_�E��e�e�d�e�g�m�[�ԜY����R�	N��E��d�d�e�d�g�m�G��H����V��^��U���u�g�d�u�i��G��H����W��^�D��d�d�e�d�f��W���Y����F�L�D��d�e�d�e�f�l�G��I����W��L����u�e�b�h�w�m�F��H����V��_�D��e�d�e�d�f�q�}���Y����[�^�D��d�e�d�e�g�l�G��I����V��B��U���g�d�u�k�u�m�F��H����V��_�D��d�d�d�e�u�}�W���K����X�^�D��e�d�e�d�g�m�G��H����W��NךU���e�d�h�u�g�l�F��I����W��_�E��e�e�d�d�{�W�W���I���F�_�D��e�d�e�d�g�l�F��I����V�d��U��g�u�k�w�g�l�F��I����W��^�D��e�d�d�w�w�}�W��K���D��_�D��d�e�d�e�g�l�G��H����D�=N��U��`�h�u�e�f�l�F��H����V��_�E��e�e�e�y�]�}�W��O���V��_�D��d�e�d�d�f�l�G��H����J�N��G��u�k�w�e�f�l�F��H����V��_�E��e�e�w�u�w�}�E��Y���V��_�E��e�d�d�d�g�m�G��H����FǻN��E��h�u�e�d�f�l�G��I����W��_�E��e�e�y�_�w�}�G��D���W��_�E��e�d�d�e�g�l�F��H���l�N�F���k�w�e�d�f�l�G��I����W��_�E��d�w�u�u�w�o�D���G����W��_�D��d�d�d�e�f�l�F��I���9F�\�F��u�e�d�d�f�m�F��H����W��_�D��d�y�_�u�w�m�C��Y����W��^�D��e�e�e�e�f�l�F��H���F�^�U��w�e�d�d�f�m�F��I����W��_�D��w�u�u�u�e�n�W���[����W��^�E��e�d�d�d�g�l�G��[��ƹF�]�H���e�d�d�d�g�l�G��I����V��^�D��y�_�u�u�g�e�J���I����W��_�D��d�d�e�e�f�m�F��U���F��W��K���e�d�d�d�g�l�F��H����V��_�D���u�u�u�g�c�}�I���I����W��_�E��d�e�d�d�g�l�F���Y���T��N��U��d�d�d�e�f�m�G��I����V��^�E���_�u�u�e�e�`�W��H����V��^�E��d�e�e�e�f�m�F��s���V��S�W��d�d�d�e�f�l�G��I����V��^�W���u�u�g�a�w�c�U��H����V��_�D��d�e�d�e�f�l�U���Y���R��
P��E��d�d�e�d�g�m�F��H����V��_�Y�ߊu�u�e�c�j�}�G��H����W��^�D��e�d�d�e�f�l�[�ԜY����Q�	N��E��d�d�e�d�f�m�F��I����V��_��U���u�g�a�u�i��G��H����W��_�E��e�d�d�e�f��W���Y����
F�L�D��d�e�d�e�g�m�G��H����W��L����u�e�e�h�w�m�F��H����V��^�E��e�d�d�e�f�q�}���Y����[�^�D��d�e�d�d�f�m�F��I����W��B��U���g�`�u�k�u�m�F��H����W��_�D��d�d�d�d�u�}�W���K����X�^�D��e�d�e�e�g�m�F��H����V��NךU���e�a�h�u�g�l�F��I����V��_�D��d�d�d�d�{�W�W���I���F�_�D��e�d�d�d�g�m�G��I����W�d��U��`�u�k�w�g�l�F��I����W��_�D��d�e�d�w�w�}�W��L���D��_�D��d�e�e�d�f�m�G��I����D�=N��U��m�h�u�e�f�l�F��H����W��^�E��d�e�d�y�]�}�W��@���V��_�D��d�d�d�d�g�m�G��I����J�N��G��u�k�w�e�f�l�F��H����W��^�D��d�e�w�u�w�}�E��Y���V��_�E��e�e�d�d�f�l�G��I����FǻN��E��h�u�e�d�f�l�G��I����W��^�E��d�d�y�_�w�}�G��D���W��_�E��d�e�e�e�f�m�F��I���l�N�C���k�w�e�d�f�l�G��H����V��^�D��e�w�u�u�w�o�A���G����W��_�D��d�e�d�e�f�m�G��I���9F�\�C��u�e�d�d�f�m�F��H����V��_�D��d�y�_�u�w�m�@��Y����W��^�D��e�d�d�d�f�l�G��I���F�^�U��w�e�d�d�f�m�F��I����W��^�E��w�u�u�u�e�k�W���[����W��^�E��e�d�d�e�f�l�G��[��ƹF�Y�H���e�d�d�d�g�l�G��H����W��^�D��y�_�u�u�g�l�J���I����W��_�D��e�d�e�d�f�m�G��U���F�� \��K���e�d�d�d�g�l�F��I����W��_�D���u�u�u�g�`�}�I���I����W��_�D��d�d�d�e�g�l�F���Y���T��N��U��d�d�d�e�f�m�F��I����W��^�D���_�u�u�e�b�`�W��H����V��^�E��e�e�e�d�g�m�G��s���V��S�W��d�d�d�e�f�l�G��H����W��_�W���u�u�g�b�w�c�U��H����V��_�E��e�e�e�d�g�l�U���Y���Q��
P��E��d�d�e�d�g�l�G��I����V��^�Y�ߊu�u�e�l�j�}�G��H����W��_�E��e�e�e�d�f�m�[�ԜY����V�	N��E��d�d�e�d�f�l�G��I����V��_��U���u�g�m�u�i��G��H����W��_�E��d�d�d�d�f��W���Y����F�L�D��d�e�d�e�f�m�G��I����W��L����u�e�f�h�w�m�F��H����V��^�E��e�d�e�e�f�q�}���Y����[�^�D��d�e�d�d�f�m�G��I����V��B��U���g�m�u�k�u�m�F��H����W��^�E��d�e�d�d�u�}�W���K����X�^�D��e�d�e�d�f�l�G��I����W��NךU���e�b�h�u�g�l�F��I����W��_�D��d�d�d�d�{�W�W���I���F�_�D��e�d�d�d�f�m�F��H����W�d��U��m�u�k�w�g�l�F��I����W��_�D��e�e�d�w�w�}�W��@���D��_�D��d�e�d�d�f�l�G��I����D�=N��U��d�h�u�e�f�l�F��H����W��_�E��e�e�e�y�]�}�W��K���V��_�D��d�e�e�e�g�l�G��I����J�N��G��u�k�w�e�f�l�F��H����V��_�D��d�d�w�u�w�}�E��Y���V��_�E��d�e�e�d�f�l�G��I����FǻN��E���h�u�e�d�f�l�G��H����V��^�E��d�e�y�_�w�}�G��D���W��_�E��e�e�d�d�g�m�G��H���l�N�L���k�w�e�d�f�l�G��I����V��_�E��d�w�u�u�w�o�N���G����W��_�D��e�e�d�e�g�l�F��I���9F�\�L��u�e�d�d�f�m�F��I����V��^�E��d�y�_�u�w�l�G��Y����W��^�D��e�e�d�d�f�l�G��H���F�_�U��w�e�d�d�f�m�F��I����V��^�E��w�u�u�u�e�m�W���[����W��^�D��d�d�d�d�f�m�F��[��ƹF�^�H���e�d�d�d�g�l�F��H����V��^�E��y�_�u�u�f�i�J���I����W��_�E��d�d�d�d�f�m�F��U���F��[��K���e�d�d�d�g�l�G��H����V��^�D���u�u�u�g�g�}�I���I����W��_�E��e�e�e�e�f�m�F���Y���T�� N��U��d�d�d�e�f�l�G��I����W��^�D���_�u�u�d�o�`�W��H����V��_�D��e�e�e�d�g�m�F��s���W��S�W��d�d�d�e�f�m�F��H����V��_�W���u�u�g�d�w�c�U��H����V��^�E��e�e�d�e�g�m�U���Y���W��
P��E��d�d�e�d�f�m�G��I����W��^�Y�ߊu�u�d�g�j�}�G��H����W��^�D��e�e�d�e�g�m�[�ԜY����U�	N��E��d�d�e�d�g�l�F��I����W��_��U���u�g�d�u�i��G��H����W��_�E��d�d�d�e�f��W���Y����F�L�D��d�e�d�d�g�l�G��I����V��L����u�d�c�h�w�m�F��H����W��_�E��d�e�e�d�f�q�}���Y����[�^�D��d�e�d�e�f�m�F��I����V��B��U���g�d�u�k�u�m�F��H����V��_�E��e�e�d�e�u�}�W���K����X�^�D��e�d�d�e�f�l�G��I����V��NךU���d�e�h�u�g�l�F��I����V��_�E��e�e�d�e�{�W�W���H���F�_�D��e�d�e�e�g�m�G��H����V�d��U��g�u�k�w�g�l�F��I����V��_�E��d�e�e�w�w�}�W��K���D��_�D��d�d�d�e�f�m�F��H����D�=N��U��a�h�u�e�f�l�F��H����V��^�D��d�d�d�y�]�}�W��L���V��_�D��d�e�e�d�g�m�G��H����J�N��G��u�k�w�e�f�l�F��H����W��^�E��e�e�w�u�w�}�E��Y���V��_�E��d�d�e�d�f�l�G��H����FǻN��D��h�u�e�d�f�l�G��H����W��^�E��d�e�y�_�w�}�F��D���W��_�E��e�e�e�e�f�l�F��I���l�N�F���k�w�e�d�f�l�G��I����W��_�E��e�w�u�u�w�o�D���G����W��_�D��d�d�d�e�g�m�G��I���9F�\�G��u�e�d�d�f�m�F��H����V��^�D��d�y�_�u�w�l�D��Y����W��^�D��e�d�d�e�g�m�G��H���F�_�U��w�e�d�d�f�m�F��I����V��_�E��w�u�u�u�e�n�W���[����W��^�D��d�d�e�e�f�l�F��[��ƹF�]�H���e�d�d�d�g�l�F��I����W��_�E��y�_�u�u�f�j�J���I����W��_�E��e�d�d�d�f�l�G��U���F��V��K���e�d�d�d�g�l�G��I����V��_�E���u�u�u�g�d�}�I���I����W��_�D��d�d�e�d�g�l�F���Y���T��N��U��d�d�d�e�f�l�F��I����W��^�D���_�u�u�d�f�`�W��H����V��_�D��d�e�d�d�g�m�G��s���W��S�W��d�d�d�e�f�m�F��I����V��^�W���u�u�g�a�w�c�U��H����V��^�E��d�d�e�e�f�l�U���Y���R��
P��E��d�d�e�d�f�l�F��H����W��_�Y�ߊu�u�d�`�j�}�G��H����W��_�E��e�e�d�d�f�l�[�ԜY����P�	N��E��d�d�e�d�g�l�G��I����V��_��U���u�g�a�u�i��G��H����W��_�E��d�d�e�e�g��W���Y����F�L�D��d�e�d�d�f�l�G��H����W��L����u�d�l�h�w�m�F��H����W��_�E��e�e�e�e�f�q�}���Y����[�^�D��d�e�d�e�f�l�F��H����W��B��U���g�`�u�k�u�m�F��H����W��^�E��d�e�d�d�u�}�W���K����X�^�D��e�d�d�e�g�m�G��H����V��NךU���d�f�h�u�g�l�F��I����V��_�E��d�e�d�e�{�W�W���H���F�_�D��e�d�d�e�g�l�G��H����V�d��U��`�u�k�w�g�l�F��I����V��^�D��d�e�d�w�w�}�W��L���D��_�D��d�d�e�e�g�l�F��H����D�=N��U��b�h�u�e�f�l�F��H����V��_�D��e�e�d�y�]�}�W��A���V��_�D��d�d�e�d�f�l�G��I����J�N��G���u�k�w�e�f�l�F��H����V��_�E��e�e�w�u�w�}�E��Y���V��_�E��d�e�d�d�g�m�G��I����FǻN��D��h�u�e�d�f�l�G��H����W��^�E��e�e�y�_�w�}�F��D���W��_�E��d�e�d�e�g�l�F��I���l�N�C���k�w�e�d�f�l�G��H����W��^�D��e�w�u�u�w�o�A���G����W��_�D��e�d�d�e�f�l�F��I���9F�\�@��u�e�d�d�f�m�F��I����V��_�E��e�y�_�u�w�l�A��Y����W��^�D��d�e�e�d�f�l�F��I���F�_�U��w�e�d�d�f�m�F��H����W��_�D��w�u�u�u�e�k�W���[����W��^�D��e�d�e�d�f�l�F��[��ƹF�X�H���e�d�d�d�g�l�F��I����V��_�D��y�_�u�u�f�m�J���I����W��_�D��d�e�e�d�g�l�G��U���F�� _��K���e�d�d�d�g�l�F��H����V��_�D���u�u�u�g�`�}�I���I����W��_�E��d�d�d�e�f�m�F���Y���T��N��U��d�d�d�e�f�l�G��H����V��_�E���_�u�u�d�c�`�W��H����V��_�D��e�d�d�e�f�l�G��s���W��S�W��d�d�d�e�f�l�F��H����V��_�W���u�u�g�b�w�c�U��H����V��_�D��d�d�d�d�f�m�U���Y���Q��
P��E��d�d�e�d�f�m�F��H����V��^�Y�ߊu�u�d�m�j�}�G��H����W��^�D��e�e�e�d�f�l�[�ԜY����_�	N��E��d�d�e�d�f�l�F��I����W��_��U���u�g�m�u�i��G��H����W��_�D��d�e�d�d�f��W���Y����F�L�D��d�e�d�d�f�m�G��H����V��L����u�d�g�h�w�m�F��H����W��^�D��e�e�d�d�f�q�}���Y����[�^�D��d�e�d�d�g�m�G��I����V��B��U���g�m�u�k�u�m�F��H����W��^�E��d�e�e�e�u�}�W���K����X�^�D��e�d�d�d�g�m�G��H����W��NךU���d�c�h�u�g�l�F��I����W��^�D��d�e�d�e�{�W�W���H���F�_�D��e�d�d�e�f�m�G��I����W�d��U��m�u�k�w�g�l�F��I����V��_�E��d�d�d�w�w�}�W��A���D��_�D��d�d�d�d�g�l�G��I����D�=N��U��e�h�u�e�f�l�F��H����W��_�E��d�e�d�y�]�}�W��H���V��_�D��d�d�e�e�g�m�F��H����J�N��G��u�k�w�e�f�l�F��H����V��_�E��d�d�w�u�w�}�E��Y���V��_�E��d�d�d�e�f�m�F��H����FǻN��D��h�u�e�d�f�l�G��H����V��^�E��d�d�y�_�w�}�F��D���W��_�E��d�e�d�e�f�m�F��H���l�N�L���k�w�e�d�f�l�G��H����W��_�E��d�w�u�u�w�o�N���G����W��_�D��d�e�e�d�f�l�G��H���9F�\�M��u�e�d�d�f�m�F��H����V��_�E��d�y�_�u�w�l�N��Y����W��^�D��d�e�d�e�f�l�G��H���F�\�U��w�e�d�d�f�m�F��H����V��_�D��w�u�u�u�e�m�W���[����W��^�D��e�e�e�d�f�l�G��[��ƹF�^�H���e�d�d�d�g�l�F��I����W��_�E��y�_�u�u�e�n�J���I����W��_�D��d�d�d�e�g�l�G��U���F��Z��K���e�d�d�d�g�l�F��I����V��^�E���u�u�u�g�g�}�I���I����W��_�D��e�e�e�e�f�l�G���Y���T��N��U��d�d�d�e�f�l�F��H����V��^�D���_�u�u�g�`�`�W��H����V��_�D��d�d�e�d�g�m�G��s���T��S�W��d�d�d�e�f�l�F��I����W��_�W���u�u�g�e�w�c�U��H����V��_�D��d�e�e�e�f�m�U���Y���W��
P��E��d�d�e�d�f�l�F��H����W��_�Y�ߊu�u�g�d�j�}�G��H����W��_�D��e�d�d�d�g�l�[�ԜY����T�	N��E��d�d�d�e�g�m�G��I����W��^��U���u�g�d�u�i��G��H����V��^�E��d�d�e�d�f��W���Y����F�L�D��d�e�e�e�g�m�F��H����W��L����u�g�`�h�w�m�F��H����V��^�D��d�d�e�d�g�q�}���Y����[�^�D��d�d�e�e�g�l�G��I����W��B��U���g�d�u�k�u�m�F��H����V��_�D��d�d�e�d�u�}�W���K����X�^�D��e�e�e�e�g�l�F��H����W��NךU���g�l�h�u�g�l�F��I����V��_�D��e�d�e�d�{�W�W���K���F�_�D��d�e�e�e�g�m�F��I����W�d��U��g�u�k�w�g�l�F��H����V��_�D��d�d�e�w�w�}�W��K���D��_�D��e�e�e�d�f�l�F��I����D�=N��U��f�h�u�e�f�l�F��I����W��^�E��d�e�e�y�]�}�W��M���V��_�D��e�e�e�d�f�m�G��H����J�N��G��u�k�w�e�f�l�F��I����W��^�E��e�e�w�u�w�}�E��Y���V��_�E��e�e�d�d�g�m�F��I����FǻN��G��h�u�e�d�f�l�G��I����V��_�D��e�e�y�_�w�}�E��D���W��_�D��e�d�e�d�g�m�F��H���l�N�G���k�w�e�d�f�l�F��I����V��_�D��e�w�u�u�w�o�D���G����W��_�E��e�e�d�e�f�l�F��H���9F�\�D��u�e�d�d�f�m�G��I����V��^�E��e�y�_�u�w�o�E��Y����W��^�E��d�d�d�d�g�l�G��H���F�\�U��w�e�d�d�f�l�G��H����W��_�D��w�u�u�u�e�n�W���[����W��_�E��e�d�e�e�f�m�G��[��ƹF�]�H���e�d�d�d�g�m�G��H����W��^�D��y�_�u�u�e�k�J���I����W��^�E��e�d�d�e�g�l�F��U���F��Y��K���e�d�d�d�f�m�G��I����W��^�E���u�u�u�g�d�}�I���I����W��^�E��d�e�d�d�g�l�G���Y���T��N��U��d�d�d�e�g�m�G��I����V��^�D���_�u�u�g�g�`�W��H����V��^�D��d�e�e�d�f�m�G��s���T��S�W��d�d�d�d�g�m�F��I����W��^�W���u�u�g�a�w�c�U��H����W��^�D��d�e�e�e�g�l�U���Y���R��
P��E��d�d�e�e�g�l�G��H����W��_�Y�ߊu�u�g�a�j�}�G��H����V��_�E��e�e�e�e�g�l�[�ԜY����S�	N��E��d�d�d�e�g�m�G��I����V��^��U���u�g�a�u�i��G��H����V��^�D��d�d�e�d�f��W���Y����F�L�D��d�e�e�e�f�m�G��H����W��L����u�g�m�h�w�m�F��H����V��^�D��d�e�e�e�f�q�}���Y����[�^�D��d�d�e�e�g�l�G��H����V��B��U���g�`�u�k�u�m�F��H����V��_�D��e�d�d�e�u�}�W���K����X�^�D��e�e�e�d�f�m�F��H����W��NךU���g�g�h�u�g�l�F��I����W��^�D��d�e�e�e�{�W�W���K���F�_�D��d�e�e�e�g�m�F��I����W�d��U��`�u�k�w�g�l�F��H����V��_�E��e�d�e�w�w�}�W��L���D��_�D��e�e�d�d�g�l�G��I����D�=N��U��c�h�u�e�f�l�F��I����W��_�E��e�e�d�y�]�}�W��N���V��_�D��e�e�e�d�g�l�G��H����J�N��G���u�k�w�e�f�l�F��I����W��_�D��d�d�w�u�w�}�E��Y���V��_�E��e�d�e�e�f�l�G��I����FǻN��G��h�u�e�d�f�l�G��I����V��_�D��d�e�y�_�w�}�E��D���W��_�D��e�d�e�e�f�l�G��I���l�N�C���k�w�e�d�f�l�F��I����W��_�E��d�w�u�u�w�o�A���G����W��_�E��d�e�e�e�g�m�G��H���9F�\�A��u�e�d�d�f�m�G��H����V��^�D��d�y�_�u�w�o�B��Y����W��^�E��d�d�d�e�g�m�G��H���F�\�U��w�e�d�d�f�l�G��H����V��_�D��w�u�u�u�e�k�W���[����W��_�E��d�e�e�e�g�m�G��[��ƹF�X�H���e�d�d�d�g�m�G��H����V��_�E��y�_�u�u�e�d�J���I����W��^�E��e�d�e�d�f�m�F��U���F�� ^��K���e�d�d�d�f�m�G��H����W��^�E���u�u�u�g�`�}�I���I����W��^�D��e�e�e�d�g�m�G���Y���T��N��U��d�d�d�e�g�m�F��H����V��^�E���_�u�u�g�d�`�W��H����V��^�D��d�e�e�e�g�l�G��s���T��S�W��d�d�d�d�g�l�G��I����W��^�W���u�u�g�b�w�c�U��H����W��_�E��e�d�d�e�g�l�U���Y���Q��
P��E��d�d�e�e�g�m�G��I����W��_�Y�ߊu�u�g�b�j�}�G��H����V��^�E��e�e�d�d�g�l�[�ԜY����^�	N��E��d�d�d�e�f�m�F��I����W��_��U���u�g�b�u�i��G��H����V��^�E��d�e�e�e�f��W���Y����F�L�D��d�e�e�e�g�m�F��H����V��L����u�g�d�h�w�m�F��H����V��^�D��d�d�d�d�g�q�}���Y����[�^�D��d�d�e�d�g�m�G��H����V��B��U���g�m�u�k�u�m�F��H����W��^�E��d�e�d�e�u�}�W���K����X�^�D��e�e�e�e�f�l�G��H����V��NךU���g�`�h�u�g�l�F��I����V��_�E��e�d�d�e�{�W�W���K���F�_�D��d�e�d�e�f�m�G��H����W�d��U��m�u�k�w�g�l�F��H����V��_�D��d�e�e�w�w�}�W��A���D��_�D��e�e�e�d�f�m�F��H����D�=N��U��l�h�u�e�f�l�F��I����W��^�E��e�d�e�y�]�}�W��I���V��_�D��e�d�d�e�g�l�G��H����J�N��G��u�k�w�e�f�l�F��I����V��_�E��d�e�w�u�w�}�E��Y���V��_�E��e�e�e�d�g�m�G��I����FǻN��G��h�u�e�d�f�l�G��I����W��^�E��d�e�y�_�w�}�E��D���W��_�D��d�d�d�e�f�m�G��I���l�N�L���k�w�e�d�f�l�F��H����W��^�D��d�w�u�u�w�o�N���G����W��_�E��e�e�d�e�g�m�F��I���9F�\�B��u�e�d�d�f�m�G��I����V��^�D��d�y�_�u�w�o�O��Y����W��^�E��d�e�e�d�g�m�F��H���F�\�U��w�e�d�d�f�l�G��H����W��^�E��w�u�u�u�e�m�W���[����W��_�E��d�d�e�e�g�l�F��[��ƹF�^�H���e�d�d�d�g�m�G��H����V��_�D��y�_�u�u�d�o�J���I����W��^�D��d�e�d�e�g�l�F��U���F��]��K���e�d�d�d�f�m�F��H����V��_�E���u�u�u�g�g�}�I���I����W��^�E��d�e�e�e�g�m�F���Y���T��N��U��d�d�d�e�g�m�G��H����W��^�E���_�u�u�f�a�`�W��H����V��^�E��e�e�d�d�g�m�F��s���U��S�W��d�d�d�d�g�l�G��H����W��^�W���u�u�g�e�w�c�U��H����W��_�E��e�d�d�d�f�l�U���Y��� V��
P��E��d�d�e�e�g�l�G��I����W��^�Y�ߊu�u�f�e�j�}�G��H����V��_�D��e�d�e�e�g�l�[�ԜY����W�	N��E��d�d�d�e�f�m�F��I����W��^��U���u�g�d�u�i��G��H����V��^�D��d�e�e�e�g��W���Y���� F�L�D��d�e�e�e�f�m�F��H����V��L����u�f�a�h�w�m�F��H����V��_�E��d�e�d�d�f�q�}���Y����[�^�D��d�d�e�d�g�m�F��I����V��B��U���g�d�u�k�u�m�F��H����W��^�E��d�e�d�d�u�}�W���K����X�^�D��e�e�e�d�f�l�G��H����V��NךU���f�m�h�u�g�l�F��I����W��^�E��e�e�e�e�{�W�W���J���F�_�D��d�e�d�e�f�l�G��H����V�d��U��g�u�k�w�g�l�F��H����V��^�D��d�d�d�w�w�}�W��K���D��_�D��e�e�d�d�f�m�G��H����D�=N��U��g�h�u�e�f�l�F��I����V��^�D��e�d�e�y�]�}�W��J���V��_�D��e�d�d�e�f�m�F��H����J�N��G��u�k�w�e�f�l�F��I����V��^�E��e�d�w�u�w�}�E��Y���V��_�E��e�d�e�d�g�m�G��I����FǻN��F��h�u�e�d�f�l�G��I����V��^�D��e�e�y�_�w�}�D��D���W��_�D��d�d�d�d�g�m�F��I���l�N�G���k�w�e�d�f�l�F��H����V��^�E��e�w�u�u�w�o�E���G����W��_�E��d�e�d�e�g�m�G��I���9F�\�E��u�e�d�d�f�m�G��H����V��^�E��e�y�_�u�w�n�F��Y����W��^�E��d�e�e�d�f�l�G��H���F�]�U��w�e�d�d�f�l�G��H����W��^�E��w�u�u�u�e�n�W���[����W��_�E��d�d�d�d�g�l�F��[��ƹF�]�H���e�d�d�d�g�m�G��H����W��_�E��y�_�u�u�d�h�J���I����W��^�D��d�e�d�e�g�l�G��U���F��X��K���e�d�d�d�f�m�F��H����V��^�E���u�u�u�g�d�}�I���I����W��^�D��d�d�d�e�g�l�G���Y���T��N��U��d�d�d�e�g�m�F��H����W��_�E���_�u�u�f�n�`�W��H����V��_�E��e�d�d�d�f�m�F��s���U��S�W��d�d�d�d�g�m�G��H����V��_�W���u�u�g�a�w�c�U��H����W��^�E��d�e�d�e�g�l�U���Y��� R��
P��E��d�d�e�e�f�m�G��H����W��^�Y�ߊu�u�f�f�j�}�G��H����V��^�D��d�e�e�e�f�m�[�ԜY����R�	N��E��d�d�d�e�g�m�F��I����V��^��U���u�g�a�u�i��G��H����V��^�D��d�e�d�d�f��W���Y����F�L�D��d�e�e�d�g�m�F��H����V��L����u�f�b�h�w�m�F��H����W��_�E��e�e�d�e�g�q�}���Y����[�^�D��d�d�e�e�g�m�F��I����W��B��U���g�a�u�k�u�m�F��H����V��^�D��d�d�d�d�u�}�W���K����X�^�D��e�e�d�e�f�l�F��H����V��NךU���f�d�h�u�g�l�F��I����V��^�E��e�d�d�d�{�W�W���J���F�_�D��d�e�e�e�f�l�G��I����W�d��U��`�u�k�w�g�l�F��H����V��^�E��e�d�e�w�w�}�W��L���D��_�D��e�d�e�d�f�m�F��I����D�=N��U��`�h�u�e�f�l�F��I����V��^�D��e�e�d�y�]�}�W��O���V��_�D��e�e�d�e�f�l�G��H����J�N��G���u�k�w�e�f�l�F��I����V��_�D��e�d�w�u�w�}�E��Y���V��_�E��d�e�e�d�g�l�G��I����FǻN��F��h�u�e�d�f�l�G��H����V��^�E��e�e�y�_�w�}�D��D���W��_�D��e�d�d�d�f�l�G��I���l�N�C���k�w�e�d�f�l�F��I����V��^�D��d�w�u�u�w�o�A���G����W��_�E��e�e�d�e�g�m�F��I���9F�\�F��u�e�d�d�f�m�G��I����V��_�E��e�y�_�u�w�n�C��Y����W��^�E��d�e�d�e�f�m�G��H���F�]�U��w�e�d�d�f�l�G��H����V��^�E��w�u�u�u�e�k�W���[����W��_�D��d�d�e�d�g�l�G��[��ƹF�X�H���e�d�d�d�g�m�F��H����V��^�E��y�_�u�u�d�e�J���I����W��^�E��d�d�e�d�g�l�G��U���F��W��K���e�d�d�d�f�m�G��H����V��^�E���u�u�u�g�`�}�I���I����W��^�E��d�d�d�d�f�l�F���Y���T��N��U��d�d�d�e�g�l�G��H����V��_�D���_�u�u�f�e�`�W��H����V��_�E��e�d�e�d�f�l�G��s���U��S�W��d�d�d�d�g�m�G��H����W��^�W���u�u�g�b�w�c�U��H����W��^�E��d�e�d�d�g�l�U���Y��� Q��
P��E��d�d�e�e�f�l�G��H����V��_�Y�ߊu�u�f�c�j�}�G��H����V��_�D��d�e�e�e�f�l�[�ԜY����Q�	N��E��d�d�d�e�g�m�F��I����V��_��U���u�g�b�u�i��G��H����V��^�D��d�e�e�e�g��W���Y����
F�L�D��d�e�e�d�f�m�F��H����V��L����u�f�e�h�w�m�F��H����W��_�E��e�e�d�e�f�q�}���Y����[�^�D��d�d�e�e�g�m�F��H����V��B��U���g�m�u�k�u�m�F��H����V��^�D��d�e�d�e�u�}�W���K����X�^�D��e�e�d�d�f�l�F��I����W��NךU���f�a�h�u�g�l�F��I����W��^�D��d�d�d�d�{�W�W���J���F�_�D��d�e�e�e�f�l�F��H����W�d��U��m�u�k�w�g�l�F��H����V��^�D��d�d�d�w�w�}�W��A���D��_�D��e�d�d�d�f�m�G��H����D�=N��U��m�h�u�e�f�l�F��I����V��^�E��e�d�e�y�]�}�W��@���V��_�D��e�e�d�e�f�l�G��H����J�N��G��u�k�w�e�f�l�F��I����V��^�E��e�d�w�u�w�}�E��Y���V��_�E��d�d�e�d�g�l�F��I����FǻN��F��h�u�e�d�f�l�G��H����V��^�D��e�e�y�_�w�}�D��D���W��_�D��e�d�d�d�g�l�F��I���l�N�L���k�w�e�d�f�l�F��I����V��^�E��e�w�u�u�w�o�N���G����W��_�E��d�e�d�d�f�l�G��I���9F�\�C��u�e�d�d�f�m�G��H����W��^�E��d�y�_�u�w�n�@��Y����W��^�E��d�e�e�d�g�l�G��H���F�]�U��w�e�d�d�f�l�G��H����W��^�E��w�u�u�u�e�d�W���[����W��_�D��d�d�d�e�f�l�F��[��ƹF�^�H���e�d�d�d�g�m�F��H����W��_�E��y�_�u�u�c�l�J���I����W��^�E��d�e�e�d�g�m�F��U���F��\��K���e�d�d�d�f�m�G��H����V��^�D���u�u�u�g�g�}�I���I����W��^�D��d�d�e�d�g�m�F���Y���T��N��U��d�d�d�e�g�l�F��H����W��^�D���_�u�u�a�b�`�W��H����V��_�E��e�d�d�d�f�l�G��s���R��S�W��d�d�d�d�g�l�G��H����V��^�W���u�u�g�e�w�c�U��H����W��_�E��e�d�e�e�f�l�U���Y���V��
P��E��d�d�e�e�f�m�G��I����W��^�Y�ߊu�u�a�l�j�}�G��H����V��^�D��d�e�e�d�f�l�[�ԜY����V�	N��E��d�d�d�e�f�m�F��I����V��^��U���u�g�d�u�i��G��H����V��^�D��d�d�d�e�f��W���Y����F�L�D��d�e�e�d�g�m�F��H����W��L����u�a�f�h�w�m�F��H����W��_�E��d�e�e�e�g�q�}���Y����[�^�D��d�d�e�d�g�m�F��I����W��B��U���g�d�u�k�u�m�F��H����W��^�D��e�d�e�e�u�}�W���K����X�^�D��e�e�d�e�f�l�F��I����V��NךU���a�b�h�u�g�l�F��I����V��_�D��e�d�e�d�{�W�W���M���F�_�D��d�e�d�e�f�m�F��I����V�d��U��d�u�k�w�g�l�F��H����V��_�D��d�d�d�w�w�}�W��K���D��_�D��e�d�e�d�f�l�F��I����D�=N��U��d�h�u�e�f�l�F��I����W��_�D��d�e�d�y�]�}�W��K���V��_�D��e�d�d�e�g�m�G��I����J�N��G��u�k�w�e�f�l�F��I����V��_�D��e�e�w�u�w�}�E��Y���V��_�E��d�e�e�d�g�l�F��H����FǻN��A���h�u�e�d�f�l�G��H����W��_�E��d�d�y�_�w�}�C��D���W��_�D��d�d�d�e�f�l�G��I���l�N�G���k�w�e�d�f�l�F��H����W��^�E��d�w�u�u�w�o�E���G����W��_�E��e�e�d�e�f�m�G��I���9F�\�L��u�e�d�d�f�m�G��I����V��^�E��d�y�_�u�w�i�G��Y����W��^�E��d�e�e�e�f�m�G��H���F�Z�U��w�e�d�d�f�l�G��H����V��^�D��w�u�u�u�e�n�W���[����W��_�D��d�e�d�d�g�m�G��[��ƹF�]�H���e�d�d�d�g�m�F��H����V��_�E��y�_�u�u�c�i�J���I����W��^�D��e�d�d�e�f�l�G��U���F��[��K���e�d�d�d�f�m�F��H����W��^�D���u�u�u�g�d�}�I���I����W��^�E��e�d�d�d�g�m�G���Y���T�� N��U��d�d�d�e�g�l�G��H����W��^�D���_�u�u�a�o�`�W��H����V��_�D��d�e�e�e�f�m�F��s���R��S�W��d�d�d�d�g�l�G��I����V��_�W���u�u�g�a�w�c�U��H����W��_�E��e�d�d�e�f�m�U���Y���R��
P��E��d�d�e�e�f�l�G��I����W��^�Y�ߊu�u�a�g�j�}�G��H����V��_�E��d�e�d�d�f�m�[�ԜY����U�	N��E��d�d�d�e�f�m�F��I����W��^��U���u�g�a�u�i��G��H����V��^�E��d�e�e�d�g��W���Y����F�L�D��d�e�e�d�f�m�F��I����W��L����u�a�c�h�w�m�F��H����W��^�E��d�d�d�e�g�q�}���Y����[�^�D��d�d�e�d�g�l�F��I����W��B��U���g�a�u�k�u�m�F��H����W��^�D��d�e�e�e�u�}�W���K����X�^�D��e�e�d�d�f�m�F��I����V��NךU���a�e�h�u�g�l�F��I����W��_�E��e�d�d�e�{�W�W���M���F�_�D��d�e�d�e�g�l�G��I����V�d��U��`�u�k�w�g�l�F��H����V��^�E��d�e�e�w�w�}�W��L���D��_�D��e�d�d�d�g�m�F��H����D�=N��U��a�h�u�e�f�l�F��I����W��^�E��e�e�d�y�]�}�W��L���V��_�D��e�d�e�d�f�l�F��I����J�N��G���u�k�w�e�f�l�F��I����V��_�E��e�d�w�u�w�}�E��Y���V��_�E��d�d�e�e�g�l�F��H����FǻN��A��h�u�e�d�f�l�G��H����W��^�E��d�d�y�_�w�}�C��D���W��_�D��d�d�e�d�g�m�F��I���l�N�C���k�w�e�d�f�l�F��H����W��_�D��d�w�u�u�w�o�A���G����W��_�E��d�e�e�d�g�l�F��H���9F�\�G��u�e�d�d�f�m�G��H����W��_�E��d�y�_�u�w�i�D��Y����W��^�E��d�d�e�e�f�l�G��H���F�Z�U��w�e�d�d�f�l�G��H����V��^�D��w�u�u�u�e�k�W���[����W��_�D��d�e�d�e�f�m�G��[��ƹF�X�H���e�d�d�d�g�m�F��H����W��^�D��y�_�u�u�c�j�J���I����W��^�D��e�e�d�e�f�m�G��U���F��V��K���e�d�d�d�f�m�F��I����V��_�E���u�u�u�g�a�}�I���I����W��^�D��e�e�d�d�f�m�G���Y���T��N��U��d�d�d�e�g�l�F��I����V��^�E���_�u�u�a�f�`�W��H����V��_�D��e�e�e�d�f�l�G��s���R��S�W��d�d�d�d�g�l�F��I����V��^�W���u�u�g�b�w�c�U��H����W��_�D��d�d�e�e�g�m�U���Y���Q��
P��E��d�d�e�e�g�m�G��H����W��_�Y�ߊu�u�a�`�j�}�G��H����V��^�E��e�d�e�d�g�m�[�ԜY����P�	N��E��d�d�d�d�g�m�G��I����W��_��U���u�g�b�u�i��G��H����W��^�D��e�d�e�d�f��W���Y����F�L�D��d�e�e�e�g�m�G��H����W��L����u�a�l�h�w�m�F��H����V��^�D��e�e�d�d�f�q�}���Y����[�^�D��d�d�d�e�g�l�G��I����W��B��U���g�m�u�k�u�m�F��H����V��_�E��e�e�e�d�u�}�W���K����X�^�D��e�e�e�e�f�m�G��H����V��NךU���a�f�h�u�g�l�F��I����V��^�E��d�d�e�d�{�W�W���M���F�_�D��d�d�e�e�g�l�F��I����W�d��U��m�u�k�w�g�l�F��H����V��^�E��e�e�d�w�w�}�W��A���D��_�D��e�e�e�d�f�l�G��H����D�=N��U��b�h�u�e�f�l�F��I����W��_�E��e�d�d�y�]�}�W��A���V��_�D��d�e�e�d�f�m�F��H����J�N��G��u�k�w�e�f�l�F��H����W��_�D��d�d�w�u�w�}�E��Y���V��_�E��e�e�d�d�g�l�G��I����FǻN��A��h�u�e�d�f�l�G��I����V��^�D��e�e�y�_�w�}�C��D���W��_�D��e�d�e�d�g�l�F��I���l�N�L���k�w�e�d�f�l�F��I����V��_�E��d�w�u�u�w�o�N���G����W��_�E��e�e�d�e�g�m�G��H���9F�\�@��u�e�d�d�f�m�G��I����W��_�E��d�y�_�u�w�i�A��Y����W��^�D��d�d�e�d�f�m�F��H���F�Z�U��w�e�d�d�f�l�F��H����V��^�E��w�u�u�u�e�d�W���[����W��_�E��e�d�d�d�g�l�F��[��ƹF�W�H���e�d�d�d�g�m�G��I����V��^�D��y�_�u�u�b�m�J���I����W��^�E��e�e�d�d�g�l�G��U���F��_��K���e�d�d�d�f�l�G��I����W��_�D���u�u�u�g�g�}�I���I����W��_�E��d�e�d�d�f�l�G���Y���T��N��U��d�d�d�e�g�m�G��H����V��_�D���_�u�u�`�c�`�W��H����V��^�D��e�e�e�d�g�m�G��s���S��S�W��d�d�d�d�f�m�F��I����V��^�W���u�u�g�e�w�c�U��H����W��^�D��d�e�d�e�f�l�U���Y���V��
P��E��d�d�e�e�g�m�F��H����W��_�Y�ߊu�u�`�m�j�}�G��H����V��^�D��e�e�d�d�f�m�[�ԜY����_�	N��E��d�d�d�d�g�m�G��I����W��^��U���u�g�d�u�i��G��H����W��^�E��d�e�e�e�g��W���Y����F�L�D��d�e�e�e�f�m�F��I����W��L����u�`�g�h�w�m�F��H����V��^�D��d�d�e�d�g�q�}���Y����[�^�D��d�d�d�e�g�l�G��I����W��B��U���g�d�u�k�u�m�F��H����V��_�E��e�d�e�d�u�}�W���K����X�^�D��e�e�e�d�g�m�F��H����W��NךU���`�c�h�u�g�l�F��I����W��_�D��e�d�e�e�{�W�W���L���F�_�D��d�d�e�e�f�l�G��H����W�d��U��d�u�k�w�g�l�F��H����V��^�E��d�e�e�w�w�}�W��H���D��_�D��e�e�d�d�g�m�F��H����D�=N��U���e�h�u�e�f�l�F��I����W��^�E��e�e�d�y�]�}�W��H���V��_�D��d�e�e�e�f�l�G��H����J�N��G��u�k�w�e�f�l�F��H����W��^�D��e�e�w�u�w�}�E��Y���V��_�E��e�d�d�e�g�m�G��H����FǻN��@��h�u�e�d�f�l�G��I����V��_�D��e�d�y�_�w�}�B��D���W��_�D��e�e�d�e�f�l�G��I���l�N�G���k�w�e�d�f�l�F��I����W��_�E��e�w�u�u�w�o�E���G����W��_�E��d�e�e�d�f�m�G��I���9F�\�M��u�e�d�d�f�m�G��H����W��^�E��d�y�_�u�w�h�N��Y����W��^�D��d�e�e�d�g�m�G��I���F�[�U��w�e�d�d�f�l�F��H����W��^�E��w�u�u�u�e�n�W���[����W��_�E��e�e�e�d�f�l�G��[��ƹF�]�H���e�d�d�d�g�m�G��I����V��^�E��y�_�u�u�b�n�J���I����W��^�E��d�d�d�d�f�m�F��U���F��Z��K���e�d�d�d�f�l�G��H����W��_�E���u�u�u�g�d�}�I���I����W��_�D��d�d�d�d�g�l�F���Y���T��N��U��d�d�d�e�g�m�F��I����W��^�D���_�u�u�`�`�`�W��H����V��^�D��d�d�d�d�g�l�G��s���S��S�W��d�d�d�d�f�m�F��I����V��^�W���u�u�g�f�w�c�U��H����W��^�D��e�e�e�d�g�m�U���Y���R��
P��E��d�d�e�e�g�l�F��I����V��^�Y�ߊu�u�`�d�j�}�G��H����V��_�D��e�e�d�d�f�m�[�ԜY����T�	N��E��d�d�d�d�g�l�F��H����W��^��U���u�g�a�u�i��G��H����W��_�D��e�d�d�d�f��W���Y����F�L�D��d�e�e�e�f�l�F��H����V��L����u�`�`�h�w�m�F��H����V��^�E��e�d�d�e�f�q�}���Y����[�^�D��d�d�d�d�g�m�F��I����W��B��U���g�a�u�k�u�m�F��H����W��^�E��d�d�d�d�u�}�W���K����X�^�D��e�e�e�e�g�l�G��I����W��NךU���`�l�h�u�g�l�F��I����V��^�E��e�d�d�d�{�W�W���L���F�_�D��d�d�d�e�f�m�F��I����V�d��U��`�u�k�w�g�l�F��H����V��_�E��d�e�d�w�w�}�W��L���D��_�D��e�e�e�e�f�l�F��H����D�=N��U���f�h�u�e�f�l�F��I����V��_�D��e�e�d�y�]�}�W��M���V��_�D��d�d�e�e�g�l�F��I����J�N��G���u�k�w�e�f�l�F��H����V��_�E��e�d�w�u�w�}�E��Y���V��_�E��e�e�d�d�g�l�G��I����FǻN��@��h�u�e�d�f�l�G��I����W��^�D��d�e�y�_�w�}�B��D���W��_�D��d�e�e�d�f�l�F��I���l�N�@���k�w�e�d�f�l�F��H����V��_�D��d�w�u�u�w�o�A���G����W��_�E��e�d�e�d�f�m�F��I���9F�\�D��u�e�d�d�f�m�G��I����W��^�E��d�y�_�u�w�h�E��Y����W��^�D��e�d�d�d�f�m�F��I���F�[�U��w�e�d�d�f�l�F��H����W��^�D��w�u�u�u�e�k�W���[����W��_�E��e�e�e�d�f�l�F��[��ƹF�X�H���e�d�d�d�g�m�G��I����V��_�E��y�_�u�u�b�k�J���I����W��^�D��e�e�d�e�f�l�F��U���F��Y��K���e�d�d�d�f�l�F��I����V��_�E���u�u�u�g�a�}�I���I����W��_�E��e�d�d�d�f�m�G���Y���T��N��U��d�d�d�e�g�m�G��I����W��_�D���_�u�u�`�g�`�W��H����V��^�D��e�d�e�d�g�l�G��s���S��S�W��d�d�d�d�f�l�F��H����W��_�W���u�u�g�b�w�c�U��H����W��_�D��e�d�e�d�f�m�U���Y���Q��
P��E��d�d�e�e�g�m�F��I����V��^�Y�ߊu�u�`�a�j�}�G��H����V��^�E��d�d�d�e�g�l�[�ԜY����S�	N��E��d�d�d�d�f�l�G��I����W��^��U���u�g�b�u�i��G��H����W��_�D��e�d�e�e�f��W���Y����F�L�D��d�e�e�e�g�l�G��H����V��L����u�`�m�h�w�m�F��H����V��_�D��d�e�d�e�g�q�}���Y����[�^�D��d�d�d�d�f�l�G��H����V��B��U���g�m�u�k�u�m�F��H����W��_�E��d�e�d�e�u�}�W���K����X�^�D��e�e�e�e�f�l�F��H����V��NךU���`�g�h�u�g�l�F��I����W��^�D��d�d�e�e�{�W�W���L���F�_�D��d�d�d�e�g�l�G��I����V�d��U��m�u�k�w�g�l�F��H����V��^�D��d�d�d�w�w�}�W��A���D��_�D��e�e�d�e�f�m�G��I����D�=N��U���c�h�u�e�f�l�F��I����V��^�D��e�d�e�y�]�}�W��N���V��_�D��d�d�e�d�f�m�F��I����J�N��G��u�k�w�e�f�l�F��H����W��_�E��e�d�w�u�w�}�E��Y���V��_�E��e�d�e�d�f�m�F��H����FǻN��@��h�u�e�d�f�l�G��I����W��_�D��e�e�y�_�w�}�B��D���W��_�D��d�e�e�e�g�m�G��H���l�N�L���k�w�e�d�f�l�F��H����W��_�D��e�w�u�u�w�o�N���G����W��_�E��d�d�d�e�f�l�G��I���9F�\�A��u�e�d�d�f�m�G��H����V��^�E��e�y�_�u�w�h�B��Y����W��^�D��e�e�d�d�g�l�F��H���F�[�U��w�e�d�d�f�l�F��I����W��^�E��w�u�u�u�e�d�W���[����W��_�E��d�e�d�d�g�m�G��[��ƹF�W�H���e�d�d�d�g�m�G��H����W��_�E��y�_�u�u�b�d�J���I����W��^�D��d�d�d�d�g�m�G��U���F��^��K���e�d�d�d�f�l�F��I����W��^�E���u�u�u�g�g�}�I���I����W��_�D��e�e�e�d�f�l�F���Y���T��N��U��d�d�d�e�g�m�F��I����W��_�E���_�u�u�c�d�`�W��H����V��^�D��e�d�e�e�g�m�G��s���P��S�W��d�d�d�d�f�l�F��H����W��_�W���u�u�g�e�w�c�U��H����W��_�E��e�d�e�d�g�l�U���Y���V��
P��E��d�d�e�e�g�l�G��I����W��_�Y�ߊu�u�c�b�j�}�G��H����V��_�D��e�e�e�d�g�l�[�ԜY����^�	N��E��d�d�d�d�f�l�F��I����V��^��U���u�g�e�u�i��G��H����W��_�D��e�d�d�d�g��W���Y����F�L�D��d�e�e�e�f�l�G��H����W��L����u�c�d�h�w�m�F��H����V��_�D��e�d�d�d�f�q�}���Y����[�^�D��d�d�d�d�f�m�G��I����V��B��U���g�d�u�k�u�m�F��H����W��^�E��d�d�d�e�u�}�W���K����X�^�D��e�e�e�d�f�m�G��I����V��NךU���c�`�h�u�g�l�F��I����W��^�D��d�d�e�d�{�W�W���O���F�_�D��d�d�d�d�f�l�F��H����W�d��U��d�u�k�w�g�l�F��H����W��^�D��e�e�e�w�w�}�W��H���D��_�D��e�e�d�d�f�m�F��I����D�=N��U��l�h�u�e�f�l�F��I����V��^�E��d�d�e�y�]�}�W��I���V��_�D��d�e�e�e�f�m�G��H����J�N��G��u�k�w�e�f�l�F��H����V��_�D��e�d�w�u�w�}�E��Y���V��_�E��d�e�e�d�f�m�G��H����FǻN��C��h�u�e�d�f�l�G��H����W��_�D��e�e�y�_�w�}�A��D���W��_�D��e�e�d�e�g�m�F��I���l�N�G���k�w�e�d�f�l�F��I����W��_�E��e�w�u�u�w�o�E���G����W��_�E��e�e�d�e�f�m�F��H���9F�\�B��u�e�d�d�f�m�G��I����V��_�E��e�y�_�u�w�k�O��Y����W��^�D��e�d�d�d�g�m�G��H���F�X�U��w�e�d�d�f�l�F��I����V��_�E��w�u�u�u�e�n�W���[����W��_�D��d�e�d�e�f�m�F��[��ƹF�]�H���e�d�d�d�g�m�F��H����W��_�D��y�_�u�u�a�o�J���I����W��^�E��e�d�e�d�g�m�G��U���F��]��K���e�d�d�d�f�l�G��H����W��^�D���u�u�u�g�d�}�I���I����W��_�E��e�d�d�e�f�m�G���Y���T��N��U��d�d�d�e�g�l�G��I����W��_�E���_�u�u�c�a�`�W��H����V��_�E��e�e�d�e�f�l�G��s���P��S�W��d�d�d�d�f�m�G��H����W��_�W���u�u�g�f�w�c�U��H����W��^�E��e�d�d�e�g�m�U���Y���U��
P��E��d�d�e�e�f�m�G��I����V��^�Y�ߊu�u�c�e�j�}�G��H����V��^�E��d�e�d�e�g�m�[�ԜY����W�	N��E��d�d�d�d�g�l�G��I����W��^��U���u�g�a�u�i��G��H����W��_�D��e�e�e�d�g��W���Y���� F�L�D��d�e�e�d�g�m�G��H����V��L����u�c�a�h�w�m�F��H����W��^�D��d�e�d�d�g�q�}���Y����[�^�D��d�d�d�e�f�l�G��I����W��B��U���g�a�u�k�u�m�F��H����V��_�D��e�d�d�e�u�}�W���K����X�^�D��e�e�d�e�g�l�F��I����V��NךU���c�m�h�u�g�l�F��I����V��^�E��e�e�d�d�{�W�W���O���F�_�D��d�d�e�d�g�l�F��H����V�d��U��`�u�k�w�g�l�F��H����W��^�D��d�d�e�w�w�}�W��L���D��_�D��e�d�e�d�f�m�G��H����D�=N��U��g�h�u�e�f�l�F��I����W��_�D��d�d�e�y�]�}�W��J���V��_�D��d�e�d�d�g�m�G��H����J�N��G���u�k�w�e�f�l�F��H����W��^�E��e�d�w�u�w�}�E��Y���V��_�E��d�e�d�d�g�m�G��H����FǻN��C��h�u�e�d�f�l�G��H����W��_�D��e�e�y�_�w�}�A��D���W��_�D��e�d�d�d�f�l�G��I���l�N�@���k�w�e�d�f�l�F��I����V��^�E��e�w�u�u�w�o�B���G����W��_�E��d�e�e�d�g�l�F��H���9F�\�E��u�e�d�d�f�m�G��H����V��^�D��e�y�_�u�w�k�F��Y����W��^�D��e�e�d�d�g�m�F��I���F�X�U��w�e�d�d�f�l�F��I����V��_�D��w�u�u�u�e�k�W���[����W��_�D��e�e�d�d�f�m�G��[��ƹF�X�H���e�d�d�d�g�m�F��I����W��_�E��y�_�u�u�a�h�J���I����W��^�E��d�e�e�e�g�l�F��U���F��X��K���e�d�d�d�f�l�G��H����W��_�E���u�u�u�g�a�}�I���I����W��_�D��e�e�d�d�f�m�F���Y���T��N��U��d�d�d�e�g�l�F��I����V��_�D���_�u�u�c�n�`�W��H����V��_�E��d�d�d�e�f�l�G��s���P��S�W��d�d�d�d�f�m�G��I����V��^�W���u�u�g�b�w�c�U��H����W��^�D��e�d�e�e�g�m�U���Y���Q��
P��E��d�d�e�e�f�l�F��I����V��^�Y�ߊu�u�c�f�j�}�G��H����V��_�D��e�d�d�d�f�m�[�ԜY����R�	N��E��d�d�d�d�g�m�F��H����V��_��U���u�g�b�u�i��G��H����W��^�D��d�e�d�d�f��W���Y����F�L�D��d�e�e�d�f�l�F��I����V��L����u�c�b�h�w�m�F��H����W��^�E��d�d�d�e�f�q�}���Y����[�^�D��d�d�d�e�f�m�F��I����V��B��U���g�b�u�k�u�m�F��H����V��^�D��e�d�d�d�u�}�W���K����X�^�D��e�e�d�d�g�l�F��I����V��NךU���c�d�h�u�g�l�F��I����W��_�E��d�d�d�e�{�W�W���O���F�_�D��d�d�e�d�f�m�F��H����V�d��U��m�u�k�w�g�l�F��H����W��_�D��d�e�e�w�w�}�W��A���D��_�D��e�d�d�e�f�m�G��I����D�=N��U��`�h�u�e�f�l�F��I����V��_�D��e�d�d�y�]�}�W��O���V��_�D��d�e�d�d�f�m�G��H����J�N��G��u�k�w�e�f�l�F��H����V��_�E��d�e�w�u�w�}�E��Y���V��_�E��d�d�d�e�g�m�G��H����FǻN��C��h�u�e�d�f�l�G��H����W��^�E��d�d�y�_�w�}�A��D���W��_�D��e�d�e�e�f�l�F��H���l�N�L���k�w�e�d�f�l�F��I����W��^�E��e�w�u�u�w�o�N���G����W��_�E��d�d�e�e�f�l�F��I���9F�\�F��u�e�d�d�f�m�G��H����V��_�D��e�y�_�u�w�k�C��Y����W��^�D��d�d�e�e�f�l�F��I���F�X�U��w�e�d�d�f�l�F��H����W��_�D��w�u�u�u�e�d�W���[����W��_�D��d�d�d�d�g�l�G��[��ƹF�W�H���e�d�d�d�g�m�F��I����V��^�D��y�_�u�u�a�e�J���I����W��^�D��e�d�d�e�f�m�F��U���F��W��K���e�d�d�d�f�l�F��I����W��_�D���u�u�u�g�g�}�I���I����W��_�E��d�d�d�d�g�l�F���Y���T��N��U��d�d�d�e�g�l�G��H����V��^�E���_�u�u�b�e�`�W��H����V��_�E��e�e�e�e�g�l�F��s���Q��S�W��d�d�d�d�f�l�G��H����W��_�W���u�u�g�e�w�c�U��H����W��_�E��e�e�d�e�g�l�U���Y���V��
P��E��d�d�e�e�f�m�G��H����V��_�Y�ߊu�u�b�c�j�}�G��H����V��^�D��e�d�d�d�f�m�[�ԜY����Q�	N��E��d�d�d�d�f�m�G��I����W��^��U���u�g�e�u�i��G��H����W��^�E��e�d�e�d�g��W���Y����
F�L�D��d�e�e�d�g�l�F��I����W��L����u�b�e�h�w�m�F��H����W��_�E��e�d�d�e�f�q�}���Y����[�^�D��d�d�d�d�g�m�F��H����W��B��U���g�d�u�k�u�m�F��H����W��_�E��d�e�e�e�u�}�W���K����X�^�D��e�e�d�e�f�m�G��H����V��NךU���b�a�h�u�g�l�F��I����V��_�E��e�d�d�e�{�W�W���N���F�_�D��d�d�d�e�f�m�F��H����V�d��U��d�u�k�w�g�l�F��H����V��_�D��d�e�d�w�w�}�W��H���D��_�D��e�d�e�e�g�m�F��I����D�=N��U��m�h�u�e�f�l�F��I����V��^�D��d�d�d�y�]�}�W��@���V��_�D��d�d�d�e�g�m�G��I����J�N��G��u�k�w�e�f�l�F��H����V��_�E��e�d�w�u�w�}�E��Y���V��_�E��d�e�e�d�f�m�F��H����FǻN��B��h�u�e�d�f�l�G��H����V��_�E��d�e�y�_�w�}�@��D���W��_�D��d�d�d�d�g�l�F��I���l�N�G���k�w�e�d�f�l�F��H����W��_�D��e�w�u�u�w�o�E���G����W��_�E��e�e�d�d�g�m�F��H���9F�\�C��u�e�d�d�f�m�G��I����W��^�D��d�y�_�u�w�j�@��Y����W��^�D��d�e�e�d�f�m�F��H���F�Y�U��w�e�d�d�f�l�F��H����V��_�D��w�u�u�u�e�o�W���[����W��_�D��d�e�d�d�f�l�G��[��ƹF� ]�H���e�d�d�d�g�m�F��H����W��_�D��y�_�u�u�`�l�J���I����W��^�D��e�d�e�e�g�m�F��U���F��\��K���e�d�d�d�f�l�F��H����V��_�D���u�u�u�g�d�}�I���I����W��_�E��e�e�e�e�f�m�G���Y���T��N��U��d�d�d�e�g�l�G��I����W��_�D���_�u�u�b�b�`�W��H����V��_�D��e�e�e�e�f�l�F��s���Q��S�W��d�d�d�d�f�l�F��H����V��_�W���u�u�g�f�w�c�U��H����W��_�E��e�d�e�e�g�l�U���Y���U��
P��E��d�d�e�e�f�l�G��H����V��^�Y�ߊu�u�b�l�j�}�G��H����V��_�E��d�e�d�e�f�l�[�ԜY����V�	N��E��d�d�d�d�f�m�G��I����V��_��U���u�g�a�u�i��G��H����W��^�D��e�e�d�d�f��W���Y����F�L�D��d�e�e�d�f�m�G��I����W��L����u�b�f�h�w�m�F��H����W��^�E��e�e�d�e�f�q�}���Y����[�^�D��d�d�d�d�g�l�F��I����W��B��U���g�a�u�k�u�m�F��H����W��_�E��e�e�d�d�u�}�W���K����X�^�D��e�e�d�d�g�l�G��H����W��NךU���b�b�h�u�g�l�F��I����W��_�D��d�d�e�e�{�W�W���N���F�_�D��d�d�d�e�g�m�F��H����W�d��U��a�u�k�w�g�l�F��H����V��_�E��e�e�d�w�w�}�W��L���D��_�D��e�d�d�d�f�m�G��H����D�=N��U��d�h�u�e�f�l�F��I����W��^�D��e�e�d�y�]�}�W��K���V��_�D��d�d�e�e�f�l�G��I����J�N��G���u�k�w�e�f�l�F��H����W��^�E��d�e�w�u�w�}�E��Y���V��_�E��d�d�d�e�g�l�F��H����FǻN��B���h�u�e�d�f�l�G��H����W��_�E��d�e�y�_�w�}�@��D���W��_�D��d�e�d�e�f�l�G��I���l�N�@���k�w�e�d�f�l�F��H����W��_�E��d�w�u�u�w�o�B���G����W��_�E��d�e�e�d�g�m�F��H���9F�\�L��u�e�d�d�f�m�G��H����V��_�E��e�y�_�u�w�j�G��Y����W��^�D��d�e�e�e�g�l�F��H���F�Y�U��w�e�d�d�f�l�F��H����W��^�D��w�u�u�u�e�k�W���[����W��_�D��e�d�d�e�g�l�F��[��ƹF� X�H���e�d�d�d�g�m�F��I����V��^�E��y�_�u�u�`�i�J���I����W��^�D��d�d�e�e�g�l�G��U���F��[��K���e�d�d�d�f�l�F��H����V��_�D���u�u�u�g�a�}�I���I����W��_�D��d�d�d�d�f�m�G���Y���T�� N��U��d�d�d�e�g�l�F��H����W��^�D���_�u�u�b�o�`�W��H����V��_�D��e�e�d�e�g�l�F��s���Q��S�W��d�d�d�d�f�l�F��I����W��_�W���u�u�g�b�w�c�U��H����W��_�D��d�d�d�d�g�m�U���Y���Q��
P��E��d�d�e�e�f�l�F��I����W��^�Y�ߊu�u�b�g�j�}�G��H����V��_�E��d�e�e�d�g�l�[�ԜY����U�	N��E��d�d�d�d�f�l�F��I����W��_��U���u�g�b�u�i��G��H����W��_�E��e�d�e�e�f��W���Y����F�L�D��d�e�e�d�f�l�G��I����W��L����u�b�c�h�w�m�F��H����W��_�E��e�d�e�e�f�q�}���Y����[�^�D��d�d�d�d�f�l�F��H����V��B��U���g�b�u�k�u�m�F��H����W��_�D��e�e�e�e�u�}�W���K����X�^�D��e�d�e�e�g�m�F��I����W��NךU���b�e�h�u�g�l�F��I����V��^�D��e�d�d�e�{�W�W���N���F�_�D��d�e�e�e�g�m�G��I����V�d��U��m�u�k�w�g�l�F��H����V��^�E��d�e�e�w�w�}�W��A���D��_�D��d�e�e�e�f�l�F��I����D�=N��U��a�h�u�e�f�l�F��H����V��^�E��e�e�d�y�]�}�W��L���V��_�D��e�e�e�d�f�m�G��H����J�N��G��u�k�w�e�f�l�F��I����W��_�E��d�d�w�u�w�}�E��Y���V��_�E��e�e�e�d�f�l�G��I����FǻN��B��h�u�e�d�f�l�G��I����W��_�E��e�d�y�_�w�}�@��D���W��_�D��e�e�e�e�g�m�G��H���l�N�L���k�w�e�d�f�l�F��I����V��^�D��e�w�u�u�w�o�N���G����W��_�D��e�d�e�d�f�l�G��I���9F�\�G��u�e�d�d�f�m�F��I����V��_�E��d�y�_�u�w�j�D��Y����W��^�E��e�e�d�e�g�l�F��H���F�Y�U��w�e�d�d�f�l�G��I����W��_�E��w�u�u�u�e�d�W���[����W��_�E��d�e�d�d�f�l�F��[��ƹF� W�H���e�d�d�d�g�l�G��H����W��_�E��y�_�u�u�`�j�J���I����W��_�E��d�e�e�e�f�l�F��U���F��V��K���e�d�d�d�f�m�G��H����V��_�D���u�u�u�g�n�}�I���I����W��^�E��d�d�d�d�f�m�G���Y���T��N��U��d�d�d�e�f�m�G��I����W��^�E���_�u�u�m�f�`�W��H����V��^�D��d�e�e�d�g�l�F��s���^��S�W��d�d�d�d�g�m�F��H����W��_�W���u�u�g�e�w�c�U��H����W��^�E��d�d�d�e�f�l�U���Y���V��
P��E��d�d�e�d�g�m�G��I����V��^�Y�ߊu�u�m�`�j�}�G��H����W��^�D��e�e�d�e�g�l�[�ԜY����P�	N��E��d�d�d�e�g�l�F��H����W��_��U���u�g�e�u�i��G��H����V��_�E��d�d�e�d�f��W���Y����F�L�D��d�e�d�e�g�m�F��H����W��L����u�m�l�h�w�m�F��H����V��^�D��e�d�d�d�g�q�}���Y����[�^�D��d�d�e�e�f�l�F��I����V��B��U���g�d�u�k�u�m�F��H����V��^�D��e�e�e�e�u�}�W���K����X�^�D��e�d�e�e�f�m�G��I����W��NךU���m�f�h�u�g�l�F��I����V��_�E��e�e�e�d�{�W�W���A���F�_�D��d�e�e�d�g�m�F��H����W�d��U��d�u�k�w�g�l�F��H����W��_�E��d�d�d�w�w�}�W��H���D��_�D��d�e�e�d�g�m�G��I����D�=N��U��b�h�u�e�f�l�F��H����W��^�D��e�d�d�y�]�}�W��A���V��_�D��e�e�d�d�f�l�F��I����J�N��G��u�k�w�e�f�l�F��I����W��^�E��d�e�w�u�w�}�E��Y���V��_�E��e�e�d�d�g�m�F��H����FǻN��M��h�u�e�d�f�l�G��I����V��^�E��e�d�y�_�w�}�O��D���W��_�D��e�e�e�e�f�m�G��H���l�N�G���k�w�e�d�f�l�F��I����W��^�E��e�w�u�u�w�o�E���G����W��_�D��d�e�d�e�g�m�G��H���9F�\�@��u�e�d�d�f�m�F��H����W��_�E��e�y�_�u�w�e�A��Y����W��^�E��e�e�d�e�f�m�G��I���F�V�U��w�e�d�d�f�l�G��I����W��_�E��w�u�u�u�e�o�W���[����W��_�E��e�e�e�d�g�l�G��[��ƹF�\�H���e�d�d�d�g�l�G��I����W��_�D��y�_�u�u�o�m�J���I����W��_�E��d�e�e�e�g�m�G��U���F��_��K���e�d�d�d�f�m�G��H����V��_�E���u�u�u�g�d�}�I���I����W��^�D��e�e�d�e�g�m�G���Y���T��N��U��d�d�d�e�f�m�F��I����W��^�D���_�u�u�m�c�`�W��H����V��^�E��d�e�d�d�f�m�G��s���^��S�W��d�d�d�d�g�m�G��I����V��^�W���u�u�g�f�w�c�U��H����W��^�D��e�e�d�e�g�l�U���Y���U��
P��E��d�d�e�d�g�l�F��H����V��_�Y�ߊu�u�m�m�j�}�G��H����W��_�D��e�e�e�e�f�l�[�ԜY���� _�	N��E��d�d�d�e�g�m�F��I����W��_��U���u�g�a�u�i��G��H����V��^�E��d�e�d�d�f��W���Y����F�L�D��d�e�d�e�f�l�F��H����W��L����u�m�g�h�w�m�F��H����V��_�D��e�d�e�e�g�q�}���Y����[�^�D��d�d�e�e�f�m�G��I����W��B��U���g�a�u�k�u�m�F��H����V��^�D��d�d�d�e�u�}�W���K����X�^�D��e�d�e�d�g�m�F��H����W��NךU���m�c�h�u�g�l�F��I����W��_�D��e�e�d�d�{�W�W���A���F�_�D��d�e�e�d�g�l�G��H����W�d��U��a�u�k�w�g�l�F��H����W��_�E��e�d�d�w�w�}�W��M���D��_�D��d�e�d�e�g�m�F��H����D�=N��U��e�h�u�e�f�l�F��H����V��^�D��d�e�d�y�]�}�W��H���V��_�D��e�e�d�d�f�l�F��I����J�N��G���u�k�w�e�f�l�F��I����W��^�D��e�e�w�u�w�}�E��Y���V��_�E��e�d�e�d�g�l�G��H����FǻN��M��h�u�e�d�f�l�G��I����V��^�E��d�d�y�_�w�}�O��D���W��_�D��e�d�e�e�f�l�G��I���l�N�@���k�w�e�d�f�l�F��I����W��^�D��e�w�u�u�w�o�B���G����W��_�D��d�d�d�e�g�m�F��I���9F�\�M��u�e�d�d�f�m�F��H����W��_�E��d�y�_�u�w�e�N��Y����W��^�E��d�e�d�e�f�m�G��H���F�V�U��w�e�d�d�f�l�G��H����W��^�E��w�u�u�u�e�k�W���[����W��_�E��d�e�e�d�g�m�F��[��ƹF�X�H���e�d�d�d�g�l�G��H����V��^�D��y�_�u�u�o�n�J���I����W��_�E��d�e�e�d�g�m�G��U���F��Z��K���e�d�d�d�f�m�G��H����V��_�D���u�u�u�g�a�}�I���I����W��^�D��d�d�d�d�f�m�G���Y���T��N��U��d�d�d�e�f�m�G��I����V��_�E���_�u�u�m�`�`�W��H����V��^�E��d�d�e�e�f�m�F��s���^��S�W��d�d�d�d�g�l�G��I����V��^�W���u�u�g�c�w�c�U��H����W��_�E��d�e�d�e�g�l�U���Y���Q��
P��E��d�d�e�d�g�m�G��H����W��_�Y�ߊu�u�m�d�j�}�G��H����W��^�D��d�e�d�e�f�l�[�ԜY����T�	N��E��d�d�d�e�f�m�F��H����V��^��U���u�g�b�u�i��G��H����V��^�E��d�e�e�d�f��W���Y����F�L�D��d�e�d�e�g�m�F��H����V��L����u�m�`�h�w�m�F��H����V��^�D��d�e�d�d�g�q�}���Y����[�^�D��d�d�e�d�g�l�F��H����W��B��U���g�b�u�k�u�m�F��H����W��^�D��e�d�d�e�u�}�W���K����X�^�D��e�d�e�e�f�m�G��H����W��NךU���m�l�h�u�g�l�F��I����V��^�D��e�e�e�d�{�W�W���A���F�_�D��d�e�d�e�g�m�G��H����W�d��U��m�u�k�w�g�l�F��H����V��_�E��d�e�e�w�w�}�W��A���D��_�D��d�e�e�d�g�m�G��H����D�=N��U��f�h�u�e�f�l�F��H����W��_�E��d�d�d�y�]�}�W��M���V��_�D��e�d�e�d�f�l�F��H����J�N��G��u�k�w�e�f�l�F��I����W��^�D��d�e�w�u�w�}�E��Y���V��_�E��e�e�d�d�f�m�F��H����FǻN��M��h�u�e�d�f�l�G��I����W��^�E��d�d�y�_�w�}�O��D���W��_�D��d�d�e�e�f�m�F��I���l�N�M���k�w�e�d�f�l�F��H����V��_�D��d�w�u�u�w�o�N���G����W��_�D��e�e�e�d�f�l�F��H���9F�\�D��u�e�d�d�f�m�F��I����V��^�E��e�y�_�u�w�e�E��Y����W��^�E��d�e�d�e�f�l�F��I���F�V�U��w�e�d�d�f�l�G��H����W��^�E��w�u�u�u�e�d�W���[����W��_�E��e�e�e�d�f�l�G��[��ƹF�W�H���e�d�d�d�g�l�G��I����W��_�E��y�_�u�u�o�k�J���I����W��_�D��d�d�d�e�g�m�G��U���F��Y��K���e�d�d�d�f�m�F��H����W��_�E���u�u�u�g�n�}�I���I����W��^�E��d�e�e�e�g�l�F���Y���T��N��U��d�d�d�e�f�m�G��H����V��_�E���_�u�u�l�g�`�W��H����V��^�D��e�e�e�e�g�m�G��s���_��S�W��d�d�d�d�g�l�F��H����V��_�W���u�u�g�e�w�c�U��H����W��_�D��e�e�d�e�f�m�U���Y���
V��
P��E��d�d�e�d�g�m�F��H����W��_�Y�ߊu�u�l�a�j�}�G��H����W��^�E��d�d�e�d�g�m�[�ԜY����S�	N��E��d�d�d�e�f�l�F��I����V��_��U���u�g�e�u�i��G��H����V��_�E��e�e�d�d�f��W���Y����F�L�D��d�e�d�e�g�l�G��I����W��L����u�l�m�h�w�m�F��H����V��_�E��d�d�d�d�g�q�}���Y����[�^�D��d�d�e�d�f�l�G��I����W��B��U���g�d�u�k�u�m�F��H����W��_�D��e�d�e�d�u�}�W���K����X�^�D��e�d�e�d�g�m�G��H����V��NךU���l�g�h�u�g�l�F��I����W��^�D��e�e�e�e�{�W�W���@���F�_�D��d�e�d�e�g�l�G��I����W�d��U��d�u�k�w�g�l�F��H����V��^�E��e�d�d�w�w�}�W��H���D��_�D��d�e�d�e�f�m�G��I����D�=N��U��c�h�u�e�f�l�F��H����V��_�D��e�d�e�y�]�}�W��N���V��_�D��e�d�e�d�g�l�G��I����J�N��G��u�k�w�e�f�l�F��I����W��^�D��e�e�w�u�w�}�E��Y���V��_�E��e�d�e�e�f�m�G��H����FǻN��L��h�u�e�d�f�l�G��I����W��_�D��e�d�y�_�w�}�N��D���W��_�D��d�e�d�d�g�m�F��H���l�N�G���k�w�e�d�f�l�F��H����W��_�E��e�w�u�u�w�o�E���G����W��_�D��d�d�e�d�g�m�G��I���9F�\�A��u�e�d�d�f�m�F��H����V��^�D��e�y�_�u�w�d�B��Y����W��^�E��e�e�d�d�g�m�F��H���F�W�U��w�e�d�d�f�l�G��I����V��^�E��w�u�u�u�e�o�W���[����W��_�E��d�d�e�d�f�l�F��[��ƹF�\�H���e�d�d�d�g�l�G��H����W��^�D��y�_�u�u�n�d�J���I����W��_�D��d�e�e�d�g�m�F��U���F��^��K���e�d�d�d�f�m�F��H����V��^�E���u�u�u�g�d�}�I���I����W��^�D��e�d�d�e�f�l�F���Y���T��N��U��d�d�d�e�f�m�F��H����V��^�D���_�u�u�l�d�`�W��H����V��^�E��d�d�d�e�f�l�F��s���_��S�W��d�d�d�d�g�l�G��H����W��^�W���u�u�g�f�w�c�U��H����W��_�E��d�d�d�e�g�l�U���Y���
U��
P��E��d�d�e�d�g�l�G��I����V��^�Y�ߊu�u�l�b�j�}�G��H����W��_�E��e�e�d�e�g�l�[�ԜY���� ^�	N��E��d�d�d�e�f�l�G��I����W��^��U���u�g�f�u�i��G��H����V��_�D��d�e�e�e�g��W���Y����F�L�D��d�e�d�e�f�m�G��I����W��L����u�l�d�h�w�m�F��H����V��^�E��d�e�d�e�f�q�}���Y����[�^�D��d�d�e�d�f�l�F��I����W��B��U���g�a�u�k�u�m�F��H����W��_�E��e�e�d�e�u�}�W���K����X�^�D��e�d�e�d�g�l�F��H����V��NךU���l�`�h�u�g�l�F��I����W��_�D��e�d�d�d�{�W�W���@���F�_�D��d�e�d�d�g�m�G��H����W�d��U��a�u�k�w�g�l�F��H����W��^�E��e�d�d�w�w�}�W��M���D��_�D��d�e�d�d�g�m�F��I����D�=N��U��l�h�u�e�f�l�F��H����W��^�D��d�d�e�y�]�}�W��I���V��_�D��e�d�d�e�g�l�G��I����J�N��G���u�k�w�e�f�l�F��I����V��_�D��d�e�w�u�w�}�E��Y���V��_�E��e�d�d�e�g�m�F��I����FǻN��L��h�u�e�d�f�l�G��I����V��^�E��e�d�y�_�w�}�N��D���W��_�D��d�d�d�d�f�m�F��H���l�N�@���k�w�e�d�f�l�F��H����V��_�E��e�w�u�u�w�o�B���G����W��_�D��d�d�d�d�g�m�F��I���9F�\�B��u�e�d�d�f�m�F��H����V��_�E��e�y�_�u�w�d�O��Y����W��^�E��e�e�e�e�f�l�G��H���F�W�U��w�e�d�d�f�l�G��I����W��^�D��w�u�u�u�e�k�W���[����W��_�D��e�e�e�d�f�l�F��[��ƹF�X�H���e�d�d�d�g�l�F��I����V��^�E��y�_�u�u�n�o�J���I����W��_�E��e�e�e�d�f�l�G��U���F��]��K���e�d�d�d�f�m�G��I����V��^�D���u�u�u�g�a�}�I���I����W��^�E��e�e�e�e�g�m�F���Y���T��N��U��d�d�d�e�f�l�G��I����W��^�E���_�u�u�l�a�`�W��H����V��_�E��d�d�e�e�g�m�F��s���_��S�W��d�d�d�d�g�m�G��I����V��_�W���u�u�g�c�w�c�U��H����W��^�E��d�d�e�d�f�m�U���Y���
P��
P��E��d�d�e�d�f�m�G��I����V��_�Y�ߊu�u�l�e�j�}�G��H����W��^�E��e�e�d�e�f�l�[�ԜY����W�	N��E��d�d�d�e�g�m�G��I����V��_��U���u�g�b�u�i��G��H����V��^�E��e�e�e�d�g��W���Y���� F�L�D��d�e�d�d�g�l�G��H����W��L����u�l�a�h�w�m�F��H����W��_�E��e�d�e�e�f�q�}���Y����[�^�D��d�d�e�e�g�m�F��I����V��B��U���g�b�u�k�u�m�F��H����V��^�D��e�d�d�e�u�}�W���K����X�^�D��e�d�d�e�f�m�F��H����W��NךU���l�m�h�u�g�l�F��I����V��^�D��e�e�d�e�{�W�W���@���F�_�D��d�e�e�e�f�l�F��I����W�d��U��m�u�k�w�g�l�F��H����V��^�E��e�e�d�w�w�}�W��A���D��_�D��d�d�e�d�f�m�F��H����D�=N��U��g�h�u�e�f�l�F��H����W��_�D��d�d�d�y�]�}�W��J���V��_�D��e�e�d�e�g�m�G��I����J�N��G��u�k�w�e�f�l�F��I����V��^�D��d�d�w�u�w�}�E��Y���V��_�E��d�e�e�e�f�m�G��I����FǻN��L��h�u�e�d�f�l�G��H����W��_�D��d�e�y�_�w�}�N��D���W��_�D��e�d�e�d�g�l�F��H���l�N�M���k�w�e�d�f�l�F��I����W��^�D��d�w�u�u�w�o�O���G����W��_�D��e�e�e�e�f�l�G��I���9F�\�E��u�e�d�d�f�m�F��I����V��_�E��e�y�_�u�w�d�F��Y����W��^�E��d�d�d�e�f�m�F��H���F�W�U��w�e�d�d�f�l�G��H����W��^�E��w�u�u�u�e�d�W���[����W��_�D��e�d�d�d�f�l�G��[��ƹF�W�H���e�d�d�d�g�l�F��I����W��_�E��y�_�u�u�n�h�J���I����W��_�E��e�e�d�e�g�m�G��U���F��X��K���e�d�d�d�f�m�G��I����V��^�E���u�u�u�g�n�}�I���I����W��^�E��e�d�e�e�g�m�F���Y���T��N��U��d�d�d�e�f�l�G��H����V��_�D���_�u�u�l�n�`�W��H����V��_�D��e�d�d�e�g�m�F��s��� V��S�W��d�d�d�d�g�m�F��H����W��_�W���u�u�f�e�w�c�U��H����W��^�D��e�d�e�d�g�m�U���Y���V��
P��E��d�d�e�d�f�m�F��H����W��_�Y�ߊu�u�e�f�j�}�G��H����W��^�D��d�e�e�d�f�m�[�ԜY����R�	N��E��d�d�d�e�g�l�F��I����W��_��U���u�f�e�u�i��G��H����V��_�D��d�e�e�d�f��W���Y����F�L�D��d�e�d�d�g�l�F��I����V��L����u�e�b�h�w�m�F��H����W��_�D��d�d�d�d�g�q�}���Y����[�^�D��d�d�e�e�g�m�G��H����W��B��U���f�e�u�k�u�m�F��H����V��^�E��d�e�e�e�u�}�W���J����X�^�D��e�d�d�d�g�m�F��I����V��NךU���e�d�h�u�g�l�F��I����W��_�E��e�e�e�e�{�W�W���I���F�_�D��d�e�e�e�g�l�G��H����V�d��U��d�u�k�w�g�l�F��H����V��_�E��d�e�d�w�w�}�W��H���D��_�D��d�d�d�e�g�m�F��I����D�=N��U��`�h�u�e�f�l�F��H����V��^�E��d�e�e�y�]�}�W��O���V��_�D��e�e�e�d�f�m�G��H����J�N��F��u�k�w�e�f�l�F��I����W��_�D��e�e�w�u�w�}�D��Y���V��_�E��d�d�e�d�f�l�G��H����FǻN��E��h�u�e�d�f�l�G��H����W��^�E��d�e�y�_�w�}�G��D���W��_�D��e�e�e�e�g�l�G��H���l�N�G���k�w�e�d�f�l�F��I����V��_�E��d�w�u�u�w�n�E���G����W��_�D��d�d�e�e�f�m�F��I���9F�]�F��u�e�d�d�f�m�F��H����V��^�E��e�y�_�u�w�m�C��Y����W��^�E��e�e�e�e�f�l�F��H���F�^�U��w�e�d�d�f�l�G��I����W��^�E��w�u�u�u�d�o�W���[����W��_�D��d�d�d�d�f�m�F��[��ƹF�\�H���e�d�d�d�g�l�F��H����V��^�E��y�_�u�u�g�e�J���I����W��_�E��d�d�e�d�g�l�F��U���F��W��K���e�d�d�d�f�m�G��H����W��_�D���u�u�u�f�d�}�I���I����W��^�D��d�e�d�d�g�m�G���Y���U��N��U��d�d�d�e�f�l�F��H����W��^�D���_�u�u�e�e�`�W��H����V��_�E��d�e�d�e�g�l�G��s��� V��S�W��d�d�d�d�g�m�F��I����V��_�W���u�u�f�f�w�c�U��H����W��^�E��d�d�e�d�f�m�U���Y���U��
P��E��d�d�e�d�f�l�G��H����W��^�Y�ߊu�u�e�c�j�}�G��H����W��_�E��e�d�d�d�f�m�[�ԜY���� Q�	N��E��d�d�d�e�g�l�G��H����V��_��U���u�f�f�u�i��G��H����V��_�D��d�e�d�d�g��W���Y����
F�L�D��d�e�d�d�f�m�G��I����V��L����u�e�e�h�w�m�F��H����W��^�E��d�e�e�d�g�q�}���Y����[�^�D��d�d�e�e�f�l�F��I����V��B��U���f�a�u�k�u�m�F��H����V��_�D��d�e�e�e�u�}�W���J����X�^�D��e�d�d�d�g�l�F��H����W��NךU���e�a�h�u�g�l�F��I����W��_�E��e�d�d�d�{�W�W���I���F�_�D��d�e�e�d�f�l�F��H����V�d��U��a�u�k�w�g�l�F��H����W��^�D��e�d�e�w�w�}�W��M���D��_�D��d�d�d�d�g�m�G��H����D�=N��U��m�h�u�e�f�l�F��H����W��_�D��d�e�d�y�]�}�W��@���V��_�D��e�e�d�e�g�m�F��I����J�N��F���u�k�w�e�f�l�F��I����V��_�D��e�e�w�u�w�}�D��Y���V��_�E��d�d�d�d�g�l�G��H����FǻN��E��h�u�e�d�f�l�G��H����V��^�E��e�d�y�_�w�}�G��D���W��_�D��e�d�d�e�g�l�G��H���l�N�@���k�w�e�d�f�l�F��I����W��^�E��d�w�u�u�w�n�B���G����W��_�D��d�d�e�d�f�l�G��I���9F�]�C��u�e�d�d�f�m�F��H����W��^�D��e�y�_�u�w�m�@��Y����W��^�E��d�d�d�e�g�m�F��I���F�^�U��w�e�d�d�f�l�G��H����V��_�D��w�u�u�u�d�h�W���[����W��_�D��e�e�e�e�f�m�G��[��ƹF�X�H���e�d�d�d�g�l�F��I����W��^�E��y�_�u�u�g�l�J���I����W��_�D��e�d�e�d�g�m�G��U���F��\��K���e�d�d�d�f�m�F��I����V��_�D���u�u�u�f�a�}�I���I����W��^�E��d�d�e�e�f�m�F���Y���U��N��U��d�d�d�e�f�l�G��H����V��^�E���_�u�u�e�b�`�W��H����V��_�E��d�d�d�d�f�m�F��s��� V��S�W��d�d�d�d�g�l�G��I����V��^�W���u�u�f�c�w�c�U��H����W��_�E��e�d�e�d�f�l�U���Y���P��
P��E��d�d�e�d�f�m�G��H����V��^�Y�ߊu�u�e�l�j�}�G��H����W��^�D��d�e�d�d�g�m�[�ԜY����V�	N��E��d�d�d�e�f�m�F��I����W��^��U���u�f�b�u�i��G��H����V��^�D��e�d�d�d�f��W���Y����F�L�D��d�e�d�d�g�l�G��H����W��L����u�e�f�h�w�m�F��H����W��_�E��e�d�d�d�g�q�}���Y����[�^�D��d�d�e�d�g�m�F��I����W��B��U���f�b�u�k�u�m�F��H����W��^�E��e�d�d�d�u�}�W���J����X�^�D��e�d�d�e�f�l�F��H����V��NךU���e�b�h�u�g�l�F��I����V��_�E��d�d�e�d�{�W�W���I���F�_�D��d�e�d�e�g�l�F��H����V�d��U��b�u�k�w�g�l�F��H����V��^�D��d�d�d�w�w�}�W��A���D��_�D��d�d�e�d�g�m�G��I����D�=N��U��d�h�u�e�f�l�F��H����W��_�D��d�e�e�y�]�}�W��K���V��_�D��e�d�e�d�g�m�F��H����J�N��F��u�k�w�e�f�l�F��I����W��_�D��e�e�w�u�w�}�D��Y���V��_�E��d�e�d�d�g�l�G��I����FǻN��E���h�u�e�d�f�l�G��H����W��_�E��d�e�y�_�w�}�G��D���W��_�D��d�d�e�e�g�l�G��H���l�N�M���k�w�e�d�f�l�F��H����W��^�D��d�w�u�u�w�n�O���G����W��_�D��e�e�e�d�g�m�G��I���9F�]�L��u�e�d�d�f�m�F��I����V��_�D��e�y�_�u�w�m�G��Y����W��^�E��d�e�e�d�f�m�G��I���F�^�U��w�e�d�d�f�l�G��H����V��^�E��w�u�u�u�d�d�W���[����W��_�D��e�e�e�e�f�l�G��[��ƹF�W�H���e�d�d�d�g�l�F��I����W��_�E��y�_�u�u�g�i�J���I����W��_�D��d�d�d�e�f�m�F��U���F��[��K���e�d�d�d�f�m�F��H����V��_�E���u�u�u�f�n�}�I���I����W��^�E��d�e�d�d�f�m�G���Y���U�� N��U��d�d�d�e�f�l�G��H����V��_�E���_�u�u�e�o�`�W��H����V��_�D��d�e�e�d�g�l�G��s��� V��S�W��d�d�d�d�g�l�F��I����W��_�W���u�u�f�e�w�c�U��H����W��_�D��d�e�e�d�f�m�U���Y���V��
P��E��d�d�e�d�f�m�F��I����V��_�Y�ߊu�u�d�g�j�}�G��H����W��^�E��d�d�d�e�f�m�[�ԜY����U�	N��E��d�d�d�e�f�l�G��I����W��_��U���u�f�e�u�i��G��H����V��_�D��d�d�e�e�f��W���Y����F�L�D��d�e�d�d�g�l�F��H����V��L����u�d�c�h�w�m�F��H����W��_�E��d�e�d�e�f�q�}���Y����[�^�D��d�d�e�d�f�l�G��I����V��B��U���f�e�u�k�u�m�F��H����W��_�E��d�e�e�e�u�}�W���J����X�^�D��e�d�d�e�f�l�G��I����V��NךU���d�e�h�u�g�l�F��I����V��_�E��d�e�e�e�{�W�W���H���F�_�D��d�e�d�d�f�l�G��I����V�d��U��d�u�k�w�g�l�F��H����W��_�E��d�e�d�w�w�}�W��H���D��_�D��d�d�d�e�g�m�F��H����D�=N��U��a�h�u�e�f�l�F��H����V��_�D��d�e�d�y�]�}�W��L���V��_�D��e�d�e�e�f�m�G��H����J�N��F��u�k�w�e�f�l�F��I����V��^�D��d�d�w�u�w�}�D��Y���V��_�E��d�d�e�d�f�l�G��I����FǻN��D��h�u�e�d�f�l�G��H����W��^�D��e�d�y�_�w�}�F��D���W��_�D��d�e�e�d�f�l�G��H���l�N�G���k�w�e�d�f�l�F��H����V��^�D��d�w�u�u�w�n�E���G����W��_�D��d�e�e�d�f�l�F��H���9F�]�G��u�e�d�d�f�m�F��H����W��^�D��e�y�_�u�w�l�D��Y����W��^�E��e�d�e�e�g�l�G��H���F�_�U��w�e�d�d�f�l�G��I����V��_�D��w�u�u�u�d�o�W���[����W��_�D��e�d�e�e�f�m�G��[��ƹF�\�H���e�d�d�d�g�l�F��I����V��_�D��y�_�u�u�f�j�J���I����W��_�D��e�e�d�e�f�l�G��U���F��V��K���e�d�d�d�f�m�F��I����W��_�E���u�u�u�f�e�}�I���I����W��^�D��e�d�e�e�g�m�G���Y���U��N��U��d�d�d�e�f�l�F��H����V��_�D���_�u�u�d�f�`�W��H����V��_�E��e�e�d�d�g�l�F��s��� W��S�W��d�d�d�d�g�l�G��H����W��_�W���u�u�f�f�w�c�U��H����W��_�D��d�e�e�d�g�m�U���Y���U��
P��E��d�d�e�d�f�l�F��I����V��_�Y�ߊu�u�d�`�j�}�G��H����W��_�D��d�d�e�d�g�l�[�ԜY���� P�	N��E��d�d�d�e�f�m�F��I����W��^��U���u�f�f�u�i��G��H����V��^�D��e�d�d�d�g��W���Y����F�L�D��d�e�d�d�f�l�F��H����V��L����u�d�l�h�w�m�F��H����W��_�D��d�e�d�d�g�q�}���Y����[�^�D��d�d�e�d�g�l�F��I����V��B��U���f�a�u�k�u�m�F��H����W��^�E��d�d�d�d�u�}�W���J����X�^�D��e�d�d�d�g�m�F��H����W��NךU���d�f�h�u�g�l�F��I����W��^�D��e�d�d�e�{�W�W���H���F�_�D��d�e�d�d�g�m�G��I����V�d��U��a�u�k�w�g�l�F��H����W��^�E��d�d�e�w�w�}�W��M���D��_�D��d�d�d�e�f�m�F��I����D�=N��U��b�h�u�e�f�l�F��H����V��_�D��d�e�e�y�]�}�W��A���V��_�D��e�d�d�d�g�l�G��I����J�N��F��u�k�w�e�f�l�F��I����W��_�E��e�e�w�u�w�}�D��Y���V��_�E��d�d�e�e�g�l�G��H����FǻN��D��h�u�e�d�f�l�G��H����V��_�D��e�e�y�_�w�}�F��D���W��_�D��d�d�d�e�g�m�G��I���l�N�@���k�w�e�d�f�l�F��H����W��_�E��e�w�u�u�w�n�B���G����W��_�D��d�e�d�d�g�l�F��I���9F�]�@��u�e�d�d�f�m�F��H����V��_�D��d�y�_�u�w�l�A��Y����W��^�E��d�e�e�e�f�m�F��I���F�_�U��w�e�d�d�f�l�G��H����W��^�E��w�u�u�u�d�h�W���[����W��_�D��d�e�d�e�g�l�F��[��ƹF�[�H���e�d�d�d�g�l�F��H����W��^�D��y�_�u�u�f�m�J���I����W��_�D��e�e�d�d�g�l�G��U���F��_��K���e�d�d�d�f�m�F��I����W��^�D���u�u�u�f�a�}�I���I����W��^�D��e�e�e�d�f�l�F���Y���U��N��U��d�d�d�e�f�l�F��I����W��_�E���_�u�u�d�c�`�W��H����V��_�D��d�e�e�d�f�m�G��s��� W��S�W��d�d�d�d�g�l�F��H����V��_�W���u�u�f�c�w�c�U��H����W��_�D��e�d�d�d�f�l�U���Y���P��
P��E��d�d�e�d�f�l�F��H����W��^�Y�ߊu�u�d�m�j�}�G��H����W��_�D��d�d�d�d�g�l�[�ԜY����_�	N��E��d�d�d�e�f�l�F��H����W��^��U���u�f�b�u�i��G��H����W��^�E��d�d�d�e�f��W���Y����F�L�D��d�e�d�e�g�m�G��H����W��L����u�d�g�h�w�m�F��H����V��^�D��e�d�e�d�f�q�}���Y����[�^�D��d�d�d�e�g�m�G��H����W��B��U���f�b�u�k�u�m�F��H����V��^�D��d�e�e�e�u�}�W���J����X�^�D��e�d�e�e�g�l�G��H����W��NךU���d�c�h�u�g�l�F��I����V��_�E��e�d�d�d�{�W�W���H���F�_�D��d�d�e�e�f�m�G��H����W�d��U��b�u�k�w�g�l�F��H����V��^�E��e�e�e�w�w�}�W��N���D��_�D��d�e�e�e�g�m�G��H����D�=N��U��e�h�u�e�f�l�F��H����V��_�D��e�e�d�y�]�}�W��H���V��_�D��d�e�e�d�g�l�G��I����J�N��F��u�k�w�e�f�l�F��H����W��_�E��d�e�w�u�w�}�D��Y���V��_�E��e�e�e�d�g�l�F��H����FǻN��D��h�u�e�d�f�l�G��I����V��^�D��d�e�y�_�w�}�F��D���W��_�D��e�e�e�e�g�l�G��I���l�N�M���k�w�e�d�f�l�F��I����W��_�E��d�w�u�u�w�n�O���G����W��_�D��e�d�e�d�f�m�F��H���9F�]�M��u�e�d�d�f�m�F��I����V��_�E��e�y�_�u�w�l�N��Y����W��^�D��e�e�e�e�f�l�F��H���F�_�U��w�e�d�d�f�l�F��I����V��_�D��w�u�u�u�d�d�W���[����W��_�E��d�d�d�e�g�l�G��[��ƹF�W�H���e�d�d�d�g�l�G��H����V��^�E��y�_�u�u�f�n�J���I����W��_�E��d�e�d�d�g�m�G��U���F��Z��K���e�d�d�d�f�l�G��H����V��_�E���u�u�u�f�n�}�I���I����W��_�E��e�d�d�d�g�m�G���Y���U��N��U��d�d�d�e�f�m�G��H����V��^�D���_�u�u�d�`�`�W��H����V��^�E��e�d�d�e�f�l�F��s��� W��S�W��d�d�d�d�f�m�G��H����V��_�W���u�u�f�l�w�c�U��H����W��^�E��e�e�d�e�f�l�U���Y���V��
P��E��d�d�e�d�g�m�G��H����V��^�Y�ߊu�u�g�d�j�}�G��H����W��^�E��e�d�d�d�f�l�[�ԜY����T�	N��E��d�d�d�d�g�l�G��I����W��_��U���u�f�e�u�i��G��H����W��_�D��d�e�d�e�g��W���Y����F�L�D��d�e�d�e�g�m�F��H����V��L����u�g�`�h�w�m�F��H����V��^�D��d�d�e�e�f�q�}���Y����[�^�D��d�d�d�e�f�m�F��H����W��B��U���f�e�u�k�u�m�F��H����V��_�E��e�e�e�e�u�}�W���J����X�^�D��e�d�e�e�g�m�F��I����W��NךU���g�l�h�u�g�l�F��I����V��^�D��d�d�d�e�{�W�W���K���F�_�D��d�d�e�d�f�l�F��I����W�d��U��d�u�k�w�g�l�F��H����W��^�E��e�d�d�w�w�}�W��H���D��_�D��d�e�e�e�f�l�G��H����D�=N��U��f�h�u�e�f�l�F��H����V��^�E��d�d�e�y�]�}�W��M���V��_�D��d�e�d�d�f�l�G��I����J�N��F��u�k�w�e�f�l�F��H����V��_�E��e�e�w�u�w�}�D��Y���V��_�E��e�e�d�e�f�l�G��I����FǻN��G��h�u�e�d�f�l�G��I����V��_�E��e�e�y�_�w�}�E��D���W��_�D��e�d�e�d�f�l�F��H���l�N�D���k�w�e�d�f�l�F��I����V��^�E��e�w�u�u�w�n�E���G����W��_�D��e�d�d�e�g�l�G��H���9F�]�D��u�e�d�d�f�m�F��I����W��_�D��e�y�_�u�w�o�E��Y����W��^�D��d�d�e�e�f�m�F��H���F�\�U��w�e�d�d�f�l�F��H����V��_�D��w�u�u�u�d�o�W���[����W��_�E��d�e�e�e�f�m�F��[��ƹF�\�H���e�d�d�d�g�l�G��H����V��^�D��y�_�u�u�e�k�J���I����W��_�E��d�e�e�e�g�l�G��U���F��Y��K���e�d�d�d�f�l�G��H����V��_�E���u�u�u�f�e�}�I���I����W��_�E��d�e�d�d�g�l�G���Y���U��N��U��d�d�d�e�f�m�G��H����W��^�D���_�u�u�g�g�`�W��H����V��^�E��e�e�e�d�f�l�G��s��� T��S�W��d�d�d�d�f�m�G��I����V��_�W���u�u�f�f�w�c�U��H����W��^�E��e�d�e�e�g�l�U���Y���U��
P��E��d�d�e�d�g�l�G��H����W��_�Y�ߊu�u�g�a�j�}�G��H����W��_�E��e�d�e�e�g�m�[�ԜY���� S�	N��E��d�d�d�d�g�m�G��I����V��_��U���u�f�f�u�i��G��H����W��^�D��d�d�d�e�g��W���Y����F�L�D��d�e�d�e�f�m�F��I����V��L����u�g�m�h�w�m�F��H����V��^�E��e�e�d�d�f�q�}���Y����[�^�D��d�d�d�e�g�l�G��I����W��B��U���f�a�u�k�u�m�F��H����V��_�E��e�d�e�e�u�}�W���J����X�^�D��e�d�e�d�g�m�F��H����V��NךU���g�g�h�u�g�l�F��I����W��_�D��e�e�e�e�{�W�W���K���F�_�D��d�d�e�e�f�m�F��I����W�d��U��a�u�k�w�g�l�F��H����V��_�E��e�e�d�w�w�}�W��M���D��_�D��d�e�d�e�f�l�G��I����D�=N��U��c�h�u�e�f�l�F��H����W��^�E��e�d�e�y�]�}�W��N���V��_�D��d�e�e�e�g�l�G��I����J�N��F��u�k�w�e�f�l�F��H����V��_�D��d�e�w�u�w�}�D��Y���V��_�E��e�d�d�e�f�m�F��H����FǻN��G��h�u�e�d�f�l�G��I����W��^�E��e�d�y�_�w�}�E��D���W��_�D��e�e�e�e�f�l�G��H���l�N�@���k�w�e�d�f�l�F��I����W��_�E��e�w�u�u�w�n�B���G����W��_�D��d�d�d�d�g�m�G��I���9F�]�A��u�e�d�d�f�m�F��H����V��_�D��e�y�_�u�w�o�B��Y����W��^�D��e�d�e�d�g�l�F��H���F�\�U��w�e�d�d�f�l�F��I����W��_�D��w�u�u�u�d�h�W���[����W��_�E��d�e�d�e�f�m�F��[��ƹF�[�H���e�d�d�d�g�l�G��H����V��^�E��y�_�u�u�e�d�J���I����W��_�E��d�e�d�e�g�l�F��U���F��^��K���e�d�d�d�f�l�G��H����V��^�E���u�u�u�f�a�}�I���I����W��_�D��d�d�e�d�g�m�F���Y���U��N��U��d�d�d�e�f�m�F��I����V��_�E���_�u�u�g�d�`�W��H����V��^�D��e�d�e�d�g�l�G��s��� T��S�W��d�d�d�d�f�m�F��H����W��_�W���u�u�f�c�w�c�U��H����W��^�E��d�e�e�d�f�m�U���Y���P��
P��E��d�d�e�d�g�l�G��I����V��_�Y�ߊu�u�g�b�j�}�G��H����W��_�E��e�d�d�e�f�m�[�ԜY����^�	N��E��d�d�d�d�g�l�G��I����W��^��U���u�f�c�u�i��G��H����W��_�D��d�d�e�e�g��W���Y����F�L�D��d�e�d�e�f�m�G��H����W��L����u�g�d�h�w�m�F��H����V��^�E��d�e�d�d�g�q�}���Y����[�^�D��d�d�d�e�f�l�F��H����W��B��U���f�b�u�k�u�m�F��H����V��_�D��d�e�d�e�u�}�W���J����X�^�D��e�d�e�d�g�l�G��H����V��NךU���g�`�h�u�g�l�F��I����W��_�E��d�d�e�e�{�W�W���K���F�_�D��d�d�e�d�f�l�G��I����W�d��U��b�u�k�w�g�l�F��H����W��_�E��d�d�d�w�w�}�W��N���D��_�D��d�e�d�d�g�m�G��I����D�=N��U��l�h�u�e�f�l�F��H����W��_�D��e�e�d�y�]�}�W��I���V��_�D��d�e�d�e�f�m�F��H����J�N��F��u�k�w�e�f�l�F��H����V��^�D��d�d�w�u�w�}�D��Y���V��_�E��e�d�d�d�g�m�F��I����FǻN��G��h�u�e�d�f�l�G��I����W��^�D��e�e�y�_�w�}�E��D���W��_�D��e�d�e�d�g�m�G��H���l�N�M���k�w�e�d�f�l�F��I����W��_�E��e�w�u�u�w�n�O���G����W��_�D��d�d�d�d�f�l�G��I���9F�]�B��u�e�d�d�f�m�F��H����V��^�E��e�y�_�u�w�o�O��Y����W��^�D��d�d�e�d�g�l�F��H���F�\�U��w�e�d�d�f�l�F��H����W��^�E��w�u�u�u�d�d�W���[����W��_�E��d�e�d�d�g�l�F��[��ƹF�W�H���e�d�d�d�g�l�G��H����V��^�D��y�_�u�u�e�o�J���I����W��_�E��d�e�d�d�f�m�F��U���F��]��K���e�d�d�d�f�l�G��H����W��^�E���u�u�u�f�n�}�I���I����W��_�D��d�d�e�d�f�l�F���Y���U��N��U��d�d�d�e�f�m�G��I����V��^�D���_�u�u�g�a�`�W��H����V��^�E��e�e�d�d�f�l�F��s��� T��S�W��d�d�d�d�f�l�G��H����W��^�W���u�u�f�l�w�c�U��H����W��_�E��d�d�e�e�g�l�U���Y���_��
P��E��d�d�e�d�g�m�G��I����V��^�Y�ߊu�u�f�e�j�}�G��H����W��^�E��e�e�e�e�f�l�[�ԜY����W�	N��E��d�d�d�d�f�m�G��I����W��_��U���u�f�e�u�i��G��H����W��^�D��e�e�d�d�f��W���Y���� F�L�D��d�e�d�e�g�m�G��I����V��L����u�f�a�h�w�m�F��H����V��^�E��e�d�e�e�f�q�}���Y����[�^�D��d�d�d�d�g�l�G��H����W��B��U���f�e�u�k�u�m�F��H����W��_�E��e�e�d�d�u�}�W���J����X�^�D��e�d�e�e�g�m�F��H����V��NךU���f�m�h�u�g�l�F��I����V��_�D��d�e�e�d�{�W�W���J���F�_�D��d�d�d�e�f�m�F��H����W�d��U��d�u�k�w�g�l�F��H����V��_�E��d�d�d�w�w�}�W��H���D��_�D��d�e�e�e�f�l�G��H����D�=N��U��g�h�u�e�f�l�F��H����W��^�E��e�e�e�y�]�}�W��J���V��_�D��d�d�e�e�g�m�F��H����J�N��F��u�k�w�e�f�l�F��H����V��^�E��e�e�w�u�w�}�D��Y���V��_�E��e�e�d�e�f�l�G��H����FǻN��F��h�u�e�d�f�l�G��I����W��^�D��d�d�y�_�w�}�D��D���W��_�D��d�e�e�e�g�l�G��I���l�N�D���k�w�e�d�f�l�F��H����W��^�D��e�w�u�u�w�n�F���G����W��_�D��e�d�d�d�g�m�G��H���9F�]�E��u�e�d�d�f�m�F��I����W��^�E��e�y�_�u�w�n�F��Y����W��^�D��e�d�e�d�g�m�F��H���F�]�U��w�e�d�d�f�l�F��I����W��^�D��w�u�u�u�d�o�W���[����W��_�E��d�e�e�e�g�l�G��[��ƹF�\�H���e�d�d�d�g�l�G��H����V��^�E��y�_�u�u�d�h�J���I����W��_�D��d�e�d�e�g�l�F��U���F��X��K���e�d�d�d�f�l�F��H����W��^�D���u�u�u�f�e�}�I���I����W��_�E��d�e�d�d�f�l�F���Y���U��N��U��d�d�d�e�f�m�G��H����V��_�D���_�u�u�f�n�`�W��H����V��^�D��e�e�d�d�f�l�F��s��� U��S�W��d�d�d�d�f�l�F��I����V��_�W���u�u�f�f�w�c�U��H����W��_�E��d�d�d�d�g�l�U���Y��� U��
P��E��d�d�e�d�g�m�G��I����W��_�Y�ߊu�u�f�f�j�}�G��H����W��^�E��d�e�d�e�g�m�[�ԜY���� R�	N��E��d�d�d�d�f�l�G��H����V��^��U���u�f�f�u�i��G��H����W��_�D��e�d�d�e�f��W���Y����F�L�D��d�e�d�e�g�m�F��I����W��L����u�f�b�h�w�m�F��H����V��^�D��d�d�d�d�g�q�}���Y����[�^�D��d�d�d�d�f�l�G��I����V��B��U���f�f�u�k�u�m�F��H����W��_�D��d�d�d�e�u�}�W���J����X�^�D��e�d�e�e�g�m�G��H����V��NךU���f�d�h�u�g�l�F��I����V��^�E��e�d�e�d�{�W�W���J���F�_�D��d�d�d�d�f�l�F��H����W�d��U��a�u�k�w�g�l�F��H����W��^�D��d�e�e�w�w�}�W��M���D��_�D��d�e�e�e�f�l�G��I����D�=N��U��`�h�u�e�f�l�F��H����V��^�E��d�d�e�y�]�}�W��O���V��_�D��d�d�d�d�f�m�F��H����J�N��F��u�k�w�e�f�l�F��H����V��^�D��d�d�w�u�w�}�D��Y���V��_�E��e�e�d�e�f�l�G��H����FǻN��F��h�u�e�d�f�l�G��I����V��^�E��d�d�y�_�w�}�D��D���W��_�D��d�d�e�d�g�m�F��I���l�N�@���k�w�e�d�f�l�F��H����W��_�D��d�w�u�u�w�n�B���G����W��_�D��e�d�d�e�f�m�F��H���9F�]�F��u�e�d�d�f�m�F��I����W��_�E��e�y�_�u�w�n�C��Y����W��^�D��d�e�d�d�g�m�F��I���F�]�U��w�e�d�d�f�l�F��H����V��^�D��w�u�u�u�d�h�W���[����W��_�E��d�e�e�d�f�l�G��[��ƹF�[�H���e�d�d�d�g�l�G��H����V��_�D��y�_�u�u�d�e�J���I����W��_�D��d�d�e�e�f�m�G��U���F��W��K���e�d�d�d�f�l�F��H����W��^�E���u�u�u�f�a�}�I���I����W��_�E��e�d�d�d�g�m�F���Y���U��N��U��d�d�d�e�f�m�G��H����W��^�D���_�u�u�f�e�`�W��H����V��^�D��e�d�e�d�g�m�G��s��� U��S�W��d�d�d�d�f�l�F��H����V��_�W���u�u�f�c�w�c�U��H����W��_�D��d�d�d�d�g�l�U���Y��� P��
P��E��d�d�e�d�g�l�G��I����W��^�Y�ߊu�u�f�c�j�}�G��H����W��_�E��e�e�e�d�f�m�[�ԜY����Q�	N��E��d�d�d�d�f�m�G��H����V��^��U���u�f�c�u�i��G��H����W��^�E��d�e�d�d�f��W���Y����
F�L�D��d�e�d�e�f�m�G��I����V��L����u�f�e�h�w�m�F��H����V��^�E��e�d�d�e�g�q�}���Y����[�^�D��d�d�d�d�g�m�G��H����W��B��U���f�b�u�k�u�m�F��H����W��^�E��e�e�d�d�u�}�W���J����X�^�D��e�d�e�d�g�l�F��H����W��NךU���f�a�h�u�g�l�F��I����W��_�D��d�d�d�e�{�W�W���J���F�_�D��d�d�d�e�f�m�F��I����W�d��U��b�u�k�w�g�l�F��H����V��^�E��e�e�d�w�w�}�W��N���D��_�D��d�e�d�e�g�m�G��H����D�=N��U��m�h�u�e�f�l�F��H����V��_�D��e�d�e�y�]�}�W��@���V��_�D��d�d�e�d�g�m�G��H����J�N��F��u�k�w�e�f�l�F��H����W��^�D��d�e�w�u�w�}�D��Y���V��_�E��e�d�e�d�f�l�F��H����FǻN��F��h�u�e�d�f�l�G��I����W��_�E��e�e�y�_�w�}�D��D���W��_�D��d�e�d�d�f�l�F��I���l�N�M���k�w�e�d�f�l�F��H����V��^�E��d�w�u�u�w�n�O���G����W��_�D��d�d�e�d�f�l�F��I���9F�]�C��u�e�d�d�f�m�F��H����V��_�E��e�y�_�u�w�n�@��Y����W��^�D��e�e�d�e�g�l�G��H���F�]�U��w�e�d�d�f�l�F��I����W��^�E��w�u�u�u�d�e�W���[����W��_�E��d�d�e�e�f�l�G��[��ƹF�W�H���e�d�d�d�g�l�G��H����V��^�E��y�_�u�u�d�l�J���I����W��_�D��e�d�e�d�f�l�G��U���F��\��K���e�d�d�d�f�l�F��I����V��^�D���u�u�u�f�n�}�I���I����W��_�D��e�e�e�d�f�l�F���Y���U��N��U��d�d�d�e�f�m�F��I����V��_�D���_�u�u�f�b�`�W��H����V��^�E��e�d�e�e�f�m�F��s��� U��S�W��d�d�d�d�f�l�G��H����W��_�W���u�u�f�l�w�c�U��H����W��_�D��d�d�e�d�f�l�U���Y��� _��
P��E��d�d�e�d�g�l�F��I����V��^�Y�ߊu�u�f�l�j�}�G��H����W��_�D��e�e�e�d�g�l�[�ԜY����V�	N��E��d�d�d�d�f�m�F��H����W��_��U���u�f�e�u�i��G��H����W��^�D��e�d�d�d�f��W���Y����F�L�D��d�e�d�e�f�l�F��I����W��L����u�a�f�h�w�m�F��H����V��^�E��d�e�d�d�g�q�}���Y����[�^�D��d�d�d�d�f�m�G��H����W��B��U���f�e�u�k�u�m�F��H����W��^�E��e�d�e�d�u�}�W���J����X�^�D��e�d�e�d�g�m�G��H����W��NךU���a�b�h�u�g�l�F��I����W��^�D��e�e�e�e�{�W�W���M���F�_�D��d�d�d�d�g�m�F��I����W�d��U��e�u�k�w�g�l�F��H����W��^�D��d�e�e�w�w�}�W��H���D��_�D��d�e�d�e�f�m�G��H����D�=N��U��d�h�u�e�f�l�F��H����V��^�D��d�d�e�y�]�}�W��K���V��_�D��d�d�d�e�f�l�G��H����J�N��F��u�k�w�e�f�l�F��H����W��_�D��d�d�w�u�w�}�D��Y���V��_�E��e�d�e�e�f�l�G��I����FǻN��A���h�u�e�d�f�l�G��I����V��^�E��d�e�y�_�w�}�C��D���W��_�D��d�d�d�d�g�m�G��I���l�N�D���k�w�e�d�f�l�F��H����W��^�D��e�w�u�u�w�n�F���G����W��_�D��d�e�d�e�g�m�F��H���9F�]�L��u�e�d�d�f�m�F��H����W��_�E��e�y�_�u�w�i�G��Y����W��^�D��d�d�d�e�g�m�F��H���F�Z�U��w�e�d�d�f�l�F��H����V��^�E��w�u�u�u�d�o�W���[����W��_�E��e�d�d�d�f�l�G��[��ƹF�\�H���e�d�d�d�g�l�G��H����V��^�D��y�_�u�u�c�i�J���I����W��_�D��e�e�e�d�f�m�F��U���F��[��K���e�d�d�d�f�l�F��I����V��^�E���u�u�u�f�e�}�I���I����W��_�D��e�d�e�d�g�m�G���Y���U�� N��U��d�d�d�e�f�m�F��I����W��^�E���_�u�u�a�o�`�W��H����V��^�D��e�d�d�d�f�m�F��s��� R��S�W��d�d�d�d�f�l�F��I����V��_�W���u�u�f�f�w�c�U��H����W��_�D��e�d�e�e�f�m�U���Y���U��
P��E��d�d�e�d�g�l�F��H����W��^�Y�ߊu�u�a�g�j�}�G��H����W��_�E��d�e�e�d�f�l�[�ԜY���� U�	N��E��d�d�d�d�f�l�F��H����V��_��U���u�f�f�u�i��G��H����W��_�E��d�e�e�d�g��W���Y����F�L�D��d�e�d�e�f�l�G��I����W��L����u�a�c�h�w�m�F��H����V��_�D��d�d�d�d�f�q�}���Y����[�^�D��d�d�d�d�f�l�F��I����V��B��U���f�f�u�k�u�m�F��H����W��_�E��d�e�d�e�u�}�W���J����X�^�D��e�d�e�d�f�l�F��H����W��NךU���a�e�h�u�g�l�F��I����W��_�E��e�d�e�e�{�W�W���M���F�_�D��d�d�d�d�f�l�F��H����W�d��U��a�u�k�w�g�l�F��H����W��_�E��e�d�d�w�w�}�W��M���D��_�D��d�d�e�e�g�m�F��I����D�=N��U��a�h�u�e�f�l�F��H����V��_�E��e�d�e�y�]�}�W��L���V��_�D��d�e�e�e�f�m�G��H����J�N��F��u�k�w�e�f�l�F��H����V��_�E��d�d�w�u�w�}�D��Y���V��_�E��d�e�e�e�f�m�F��I����FǻN��A��h�u�e�d�f�l�G��H����W��_�D��e�d�y�_�w�}�C��D���W��_�D��e�e�e�e�g�m�F��H���l�N�@���k�w�e�d�f�l�F��I����V��_�D��e�w�u�u�w�n�B���G����W��_�D��e�e�d�e�g�m�G��I���9F�]�G��u�e�d�d�f�m�F��I����W��^�D��d�y�_�u�w�i�D��Y����W��^�D��e�d�e�e�f�m�F��H���F�Z�U��w�e�d�d�f�l�F��I����W��^�D��w�u�u�u�d�h�W���[����W��_�D��e�e�d�e�f�m�F��[��ƹF�[�H���e�d�d�d�g�l�F��I����W��_�E��y�_�u�u�c�j�J���I����W��_�E��d�d�e�e�g�l�G��U���F��V��K���e�d�d�d�f�l�G��H����V��^�D���u�u�u�f�b�}�I���I����W��_�E��d�e�d�e�f�l�F���Y���U��N��U��d�d�d�e�f�l�G��H����V��^�E���_�u�u�a�f�`�W��H����V��_�E��d�e�e�d�g�m�F��s��� R��S�W��d�d�d�d�f�m�G��H����W��^�W���u�u�f�c�w�c�U��H����W��^�E��d�d�e�d�f�m�U���Y���P��
P��E��d�d�e�d�f�m�F��I����V��_�Y�ߊu�u�a�`�j�}�G��H����W��^�E��e�e�e�e�f�l�[�ԜY����P�	N��E��d�d�d�d�g�m�G��I����W��_��U���u�f�c�u�i��G��H����W��^�E��d�d�e�e�g��W���Y����F�L�D��d�e�d�d�g�l�G��I����V��L����u�a�l�h�w�m�F��H����W��_�E��e�e�d�e�f�q�}���Y����[�^�D��d�d�d�e�g�m�G��I����W��B��U���f�b�u�k�u�m�F��H����V��^�D��d�e�e�e�u�}�W���J����X�^�D��e�d�d�e�f�l�G��I����W��NךU���a�f�h�u�g�l�F��I����V��_�E��d�e�d�e�{�W�W���M���F�_�D��d�d�e�e�f�m�G��H����V�d��U��b�u�k�w�g�l�F��H����V��^�D��e�d�d�w�w�}�W��N���D��_�D��d�d�e�d�g�l�G��H����D�=N��U��b�h�u�e�f�l�F��H����W��^�E��e�d�e�y�]�}�W��A���V��_�D��d�e�e�d�f�m�G��I����J�N��F��u�k�w�e�f�l�F��H����W��_�D��e�d�w�u�w�}�D��Y���V��_�E��d�e�d�d�g�l�F��I����FǻN��A��h�u�e�d�f�l�G��H����W��^�E��d�d�y�_�w�}�C��D���W��_�D��e�e�d�e�f�l�G��H���l�N�M���k�w�e�d�f�l�F��I����W��_�D��e�w�u�u�w�n�O���G����W��_�D��e�d�d�d�f�m�G��H���9F�]�@��u�e�d�d�f�m�F��I����V��^�E��d�y�_�u�w�i�A��Y����W��^�D��d�e�e�d�g�l�F��I���F�Z�U��w�e�d�d�f�l�F��H����W��_�D��w�u�u�u�d�e�W���[����W��_�D��e�e�e�d�f�m�F��[��ƹF�V�H���e�d�d�d�g�l�F��I����V��_�D��y�_�u�u�c�m�J���I����W��_�E��e�d�d�e�g�l�G��U���F��_��K���e�d�d�d�f�l�G��I����W��_�E���u�u�u�f�n�}�I���I����W��_�E��d�d�e�d�f�l�F���Y���U��N��U��d�d�d�e�f�l�G��H����W��^�D���_�u�u�a�c�`�W��H����V��_�D��d�d�d�d�g�l�G��s��� R��S�W��d�d�d�d�f�m�F��H����V��^�W���u�u�f�l�w�c�U��H����W��^�E��e�e�d�e�g�m�U���Y���_��
P��E��d�d�e�d�f�m�G��I����W��_�Y�ߊu�u�a�m�j�}�G��H����W��^�D��d�e�e�d�g�m�[�ԜY����
_�	N��E��d�d�d�d�g�l�F��I����V��_��U���u�f�e�u�i��G��H����W��_�E��d�d�e�d�f��W���Y����F�L�D��d�e�d�d�g�m�G��I����W��L����u�`�g�h�w�m�F��H����W��^�E��e�d�d�e�f�q�}���Y����[�^�D��d�d�d�e�f�l�G��I����W��B��U���f�e�u�k�u�m�F��H����V��_�D��e�e�d�d�u�}�W���J����X�^�D��e�d�d�e�g�l�G��H����V��NךU���`�c�h�u�g�l�F��I����V��_�E��e�d�e�e�{�W�W���L���F�_�D��d�d�e�d�f�l�F��I����V�d��U��e�u�k�w�g�l�F��H����W��^�E��e�d�e�w�w�}�W��I���D��_�D��d�d�e�d�g�l�F��H����D�=N��U���e�h�u�e�f�l�F��H����W��^�E��d�d�e�y�]�}�W��H���V��_�D��d�e�d�e�f�l�F��I����J�N��F��u�k�w�e�f�l�F��H����V��^�E��e�d�w�u�w�}�D��Y���V��_�E��d�e�d�d�g�m�F��I����FǻN��@��h�u�e�d�f�l�G��H����W��_�D��e�e�y�_�w�}�B��D���W��_�D��e�d�e�e�g�l�F��H���l�N�D���k�w�e�d�f�l�F��I����W��_�E��d�w�u�u�w�n�F���G����W��_�D��e�d�d�e�f�m�G��I���9F�]�M��u�e�d�d�f�m�F��I����W��_�D��d�y�_�u�w�h�N��Y����W��^�D��d�d�e�e�g�m�F��I���F�[�U��w�e�d�d�f�l�F��H����W��^�D��w�u�u�u�d�o�W���[����W��_�D��d�e�d�e�g�m�F��[��ƹF�\�H���e�d�d�d�g�l�F��H����W��^�D��y�_�u�u�b�n�J���I����W��_�E��d�d�e�e�g�l�G��U���F��Z��K���e�d�d�d�f�l�G��H����W��_�E���u�u�u�f�e�}�I���I����W��_�E��d�e�d�e�g�l�G���Y���U��N��U��d�d�d�e�f�l�G��H����V��_�E���_�u�u�`�`�`�W��H����V��_�D��e�d�d�d�g�l�G��s��� S��S�W��d�d�d�d�f�m�F��H����W��_�W���u�u�f�g�w�c�U��H����W��^�D��d�e�d�e�f�l�U���Y���U��
P��E��d�d�e�d�f�m�F��H����W��_�Y�ߊu�u�`�d�j�}�G��H����W��_�E��e�d�e�d�f�m�[�ԜY���� T�	N��E��d�d�d�d�g�m�G��I����V��^��U���u�f�f�u�i��G��H����W��^�E��d�e�d�d�g��W���Y����F�L�D��d�e�d�d�f�m�G��H����W��L����u�`�`�h�w�m�F��H����W��^�D��d�e�e�e�g�q�}���Y����[�^�D��d�d�d�e�g�m�F��I����W��B��U���f�f�u�k�u�m�F��H����V��^�E��d�e�d�d�u�}�W���J����X�^�D��e�d�d�d�g�l�F��I����W��NךU���`�l�h�u�g�l�F��I����W��_�D��e�e�e�d�{�W�W���L���F�_�D��d�d�e�e�g�l�G��H����W�d��U��a�u�k�w�g�l�F��H����V��_�E��d�d�d�w�w�}�W��M���D��_�D��d�d�d�e�f�l�F��H����D�=N��U���f�h�u�e�f�l�F��H����V��^�D��e�d�d�y�]�}�W��M���V��_�D��d�e�e�d�g�m�F��H����J�N��F��u�k�w�e�f�l�F��H����W��_�E��e�d�w�u�w�}�D��Y���V��_�E��d�d�e�e�g�l�F��H����FǻN��@��h�u�e�d�f�l�G��H����V��^�D��d�d�y�_�w�}�B��D���W��_�D��e�e�d�d�f�m�G��H���l�N�A���k�w�e�d�f�l�F��I����V��_�E��e�w�u�u�w�n�B���G����W��_�D��d�e�d�d�g�l�G��I���9F�]�D��u�e�d�d�f�m�F��H����W��_�E��e�y�_�u�w�h�E��Y����W��^�D��e�d�d�e�f�m�G��I���F�[�U��w�e�d�d�f�l�F��I����V��^�E��w�u�u�u�d�h�W���[����W��_�D��e�d�d�e�g�l�G��[��ƹF�[�H���e�d�d�d�g�l�F��H����W��^�D��y�_�u�u�b�k�J���I����W��_�E��e�e�d�d�f�m�G��U���F��Y��K���e�d�d�d�f�l�G��I����V��^�D���u�u�u�f�b�}�I���I����W��_�D��e�e�d�e�g�m�F���Y���U��N��U��d�d�d�e�f�l�F��I����V��^�D���_�u�u�`�g�`�W��H����V��_�E��d�d�e�d�f�m�F��s��� S��S�W��d�d�d�d�f�m�G��I����W��^�W���u�u�f�c�w�c�U��H����W��^�D��e�d�d�e�g�l�U���Y���P��
P��E��d�d�e�d�f�l�F��H����W��_�Y�ߊu�u�`�a�j�}�G��H����W��_�E��e�e�d�e�g�l�[�ԜY����S�	N��E��d�d�d�d�g�m�G��H����V��_��U���u�f�c�u�i��G��H����W��^�D��d�d�d�e�g��W���Y����F�L�D��d�e�d�d�f�l�G��I����V��L����u�`�m�h�w�m�F��H����W��_�E��d�e�d�d�g�q�}���Y����[�^�D��d�d�d�e�g�l�G��I����V��B��U���f�b�u�k�u�m�F��H����V��_�D��e�d�d�e�u�}�W���J����X�^�D��e�d�d�d�f�m�G��I����V��NךU���`�g�h�u�g�l�F��I����W��^�E��e�d�e�e�{�W�W���L���F�_�D��d�d�e�e�f�l�F��I����W�d��U��b�u�k�w�g�l�F��H����V��^�D��d�d�e�w�w�}�W��N���D��_�D��d�d�d�d�f�l�G��H����D�=N��U���c�h�u�e�f�l�F��H����W��_�D��d�d�d�y�]�}�W��N���V��_�D��d�e�e�d�f�m�G��H����J�N��F��u�k�w�e�f�l�F��H����W��_�E��d�e�w�u�w�}�D��Y���V��_�E��d�d�d�d�f�m�G��H����FǻN��@��h�u�e�d�f�l�G��H����V��^�E��d�e�y�_�w�}�B��D���W��_�D��e�d�e�e�f�l�F��H���l�N�M���k�w�e�d�f�l�F��I����V��^�D��d�w�u�u�w�n�O���G����W��_�D��d�e�e�d�f�l�G��H���9F�]�A��u�e�d�d�f�m�F��H����V��_�D��e�y�_�u�w�h�B��Y����W��^�D��d�e�d�e�f�m�G��I���F�[�U��w�e�d�d�f�l�F��H����W��^�D��w�u�u�u�d�e�W���[����W��_�D��e�d�e�d�g�l�F��[��ƹF�V�H���e�d�d�d�g�l�F��I����V��^�E��y�_�u�u�b�d�J���I����W��_�E��e�e�d�d�g�m�F��U���F��^��K���e�d�d�d�f�l�G��I����W��_�D���u�u�u�f�n�}�I���I����W��_�D��d�e�d�d�g�m�F���Y���U��N��U��d�d�d�e�f�l�F��H����W��_�D���_�u�u�`�d�`�W��H����V��_�D��e�e�e�d�f�l�F��s��� S��S�W��d�d�d�d�f�m�F��I����W��_�W���u�u�f�l�w�c�U��H����W��^�E��d�d�e�e�f�l�U���Y���_��
P��E��d�d�e�d�f�l�G��H����W��_�Y�ߊu�u�`�b�j�}�G��H����W��_�D��e�d�e�d�g�m�[�ԜY����
^�	N��E��d�d�d�d�g�l�F��I����W��^��U���u�f�l�u�i��G��H����W��_�E��e�e�d�d�f��W���Y����F�L�D��d�e�d�d�f�m�F��I����W��L����u�c�d�h�w�m�F��H����W��^�E��e�e�d�e�f�q�}���Y����[�^�D��d�d�d�e�f�l�G��H����V��B��U���f�e�u�k�u�m�F��H����V��_�E��e�d�e�d�u�}�W���J����X�^�D��e�d�d�d�g�l�G��H����W��NךU���c�`�h�u�g�l�F��I����W��_�E��e�e�e�e�{�W�W���O���F�_�D��d�d�e�d�f�l�F��H����W�d��U��e�u�k�w�g�l�F��H����W��^�D��e�e�e�w�w�}�W��I���D��_�D��d�d�d�d�g�m�F��H����D�=N��U��l�h�u�e�f�l�F��H����W��_�E��d�d�e�y�]�}�W��I���V��_�D��d�e�d�e�f�m�F��I����J�N��F��u�k�w�e�f�l�F��H����V��_�D��d�d�w�u�w�}�D��Y���V��_�E��d�d�d�e�f�l�G��I����FǻN��C��h�u�e�d�f�l�G��H����V��_�D��d�d�y�_�w�}�A��D���W��_�D��e�d�e�e�g�l�G��H���l�N�D���k�w�e�d�f�l�F��I����V��^�D��d�w�u�u�w�n�F���G����W��_�D��d�d�d�d�g�l�G��I���9F�]�B��u�e�d�d�f�m�F��H����V��^�E��e�y�_�u�w�k�O��Y����W��^�D��d�e�d�d�f�l�F��I���F�X�U��w�e�d�d�f�l�F��H����V��^�D��w�u�u�u�d�o�W���[����W��_�D��d�d�d�d�g�l�G��[��ƹF�\�H���e�d�d�d�g�l�F��H����W��_�D��y�_�u�u�a�o�J���I����W��_�E��d�e�e�e�g�l�G��U���F��]��K���e�d�d�d�f�l�G��H����V��^�E���u�u�u�f�e�}�I���I����W��_�D��e�e�e�e�g�l�G���Y���U��N��U��d�d�d�e�f�l�F��I����W��^�E���_�u�u�c�a�`�W��H����V��_�D��d�e�e�d�f�l�F��s��� P��S�W��d�d�d�d�f�m�F��H����W��_�W���u�u�f�g�w�c�U��H����W��^�D��e�d�e�e�g�l�U���Y���T��
P��E��d�d�e�d�f�l�F��I����V��_�Y�ߊu�u�c�e�j�}�G��H����W��_�D��d�e�d�e�f�l�[�ԜY���� W�	N��E��d�d�d�d�g�l�F��I����W��_��U���u�f�f�u�i��G��H����W��_�D��e�e�d�e�g��W���Y���� F�L�D��d�e�d�d�f�l�F��I����V��L����u�c�a�h�w�m�F��H����W��_�D��e�e�d�e�g�q�}���Y����[�^�D��d�d�d�d�g�m�G��I����W��B��U���f�f�u�k�u�m�F��H����W��^�E��d�d�d�e�u�}�W���J����X�^�D��e�d�d�e�g�m�F��I����V��NךU���c�m�h�u�g�l�F��I����V��^�D��e�d�d�d�{�W�W���O���F�_�D��d�d�d�e�g�l�F��I����V�d��U��a�u�k�w�g�l�F��H����V��_�E��d�d�d�w�w�}�W��M���D��_�D��d�d�e�e�g�l�G��I����D�=N��U��g�h�u�e�f�l�F��H����V��^�D��d�d�e�y�]�}�W��J���V��_�D��d�d�e�e�g�l�F��I����J�N��F��u�k�w�e�f�l�F��H����V��^�D��e�e�w�u�w�}�D��Y���V��_�E��d�e�e�d�f�l�G��H����FǻN��C��h�u�e�d�f�l�G��H����W��_�E��e�d�y�_�w�}�A��D���W��_�D��d�e�e�d�f�m�F��I���l�N�A���k�w�e�d�f�l�F��H����W��_�D��e�w�u�u�w�n�C���G����W��_�D��e�e�d�d�f�m�F��H���9F�]�E��u�e�d�d�f�m�F��I����V��_�D��d�y�_�u�w�k�F��Y����W��^�D��e�d�e�e�g�m�G��H���F�X�U��w�e�d�d�f�l�F��I����W��_�E��w�u�u�u�d�h�W���[����W��_�D��e�e�e�e�f�m�G��[��ƹF�[�H���e�d�d�d�g�l�F��I����V��^�D��y�_�u�u�a�h�J���I����W��_�D��d�d�e�d�g�m�G��U���F��X��K���e�d�d�d�f�l�F��H����W��_�D���u�u�u�f�b�}�I���I����W��_�E��d�e�e�e�f�m�G���Y���U��N��U��d�d�d�e�f�l�G��H����W��^�E���_�u�u�c�n�`�W��H����V��_�E��e�e�d�d�f�m�G��s��� P��S�W��d�d�d�d�f�l�G��I����V��^�W���u�u�f�c�w�c�U��H����W��_�E��e�d�e�d�g�l�U���Y���P��
P��E��d�d�e�d�f�m�G��I����W��^�Y�ߊu�u�c�f�j�}�G��H����W��^�D��e�e�e�e�g�m�[�ԜY����R�	N��E��d�d�d�d�f�m�F��H����W��^��U���u�f�c�u�i��G��H����W��^�E��d�d�e�e�g��W���Y����F�L�D��d�e�d�d�g�l�G��H����V��L����u�c�b�h�w�m�F��H����W��_�E��d�e�d�d�g�q�}���Y����[�^�D��d�d�d�d�g�m�G��H����V��B��U���f�c�u�k�u�m�F��H����W��^�E��e�e�d�d�u�}�W���J����X�^�D��e�d�d�e�f�m�G��I����W��NךU���c�d�h�u�g�l�F��I����V��^�E��d�d�e�e�{�W�W���O���F�_�D��d�d�d�e�g�l�F��I����V�d��U��b�u�k�w�g�l�F��H����V��^�D��e�d�d�w�w�}�W��N���D��_�D��d�d�e�d�f�m�F��H����D�=N��U��`�h�u�e�f�l�F��H����W��_�D��d�d�e�y�]�}�W��O���V��_�D��d�d�e�e�g�l�F��H����J�N��F��u�k�w�e�f�l�F��H����V��^�D��e�e�w�u�w�}�D��Y���V��_�E��d�e�d�d�g�l�F��H����FǻN��C��h�u�e�d�f�l�G��H����W��_�D��e�e�y�_�w�}�A��D���W��_�D��d�e�e�d�f�l�F��I���l�N�M���k�w�e�d�f�l�F��H����V��_�E��d�w�u�u�w�n�O���G����W��_�D��e�d�e�e�f�l�G��I���9F�]�F��u�e�d�d�f�m�F��I����W��_�D��e�y�_�u�w�k�C��Y����W��^�D��e�d�e�d�f�m�G��I���F�X�U��w�e�d�d�f�l�F��I����V��^�E��w�u�u�u�d�e�W���[����W��_�D��d�e�e�d�f�m�G��[��ƹF�V�H���e�d�d�d�g�l�F��H����W��^�E��y�_�u�u�a�e�J���I����W��_�D��d�d�d�d�f�m�F��U���F��W��K���e�d�d�d�f�l�F��H����W��_�E���u�u�u�f�n�}�I���I����W��_�E��d�e�d�e�f�l�G���Y���U��N��U��d�d�d�e�f�l�G��H����V��^�D���_�u�u�c�e�`�W��H����V��_�E��e�d�d�e�g�m�F��s��� P��S�W��d�d�d�d�f�l�G��H����W��^�W���u�u�f�l�w�c�U��H����W��_�D��e�d�d�e�g�m�U���Y���_��
P��E��d�d�e�d�f�m�F��H����V��_�Y�ߊu�u�c�c�j�}�G��H����W��^�D��d�e�d�d�g�l�[�ԜY����
Q�	N��E��d�d�d�d�f�l�G��I����V��_��U���u�f�l�u�i��G��H����W��_�E��d�e�e�d�g��W���Y����
F�L�D��d�e�d�d�g�m�G��I����W��L����u�b�e�h�w�m�F��H����W��^�E��d�e�d�d�g�q�}���Y����[�^�D��d�d�d�d�f�m�F��H����V��B��U���f�e�u�k�u�m�F��H����W��^�E��e�e�e�e�u�}�W���J����X�^�D��e�d�d�e�g�m�F��I����V��NךU���b�a�h�u�g�l�F��I����V��^�D��d�d�d�d�{�W�W���N���F�_�D��d�d�d�d�g�m�G��I����V�d��U��e�u�k�w�g�l�F��H����W��^�E��d�e�e�w�w�}�W��I���D��_�D��d�d�e�e�f�l�G��I����D�=N��U��m�h�u�e�f�l�F��H����V��_�D��d�e�e�y�]�}�W��@���V��_�D��d�d�d�e�g�l�F��H����J�N��F��u�k�w�e�f�l�F��H����V��^�E��e�d�w�u�w�}�D��Y���V��_�E��d�e�e�d�g�l�F��H����FǻN��B��h�u�e�d�f�l�G��H����W��_�E��d�e�y�_�w�}�@��D���W��_�D��d�d�e�d�f�m�F��I���l�N�D���k�w�e�d�f�l�F��H����V��^�E��d�w�u�u�w�n�F���G����W��_�D��e�e�e�e�g�l�F��I���9F�]�C��u�e�d�d�f�m�F��I����W��^�D��d�y�_�u�w�j�@��Y����W��^�D��d�d�e�d�g�l�F��I���F�Y�U��w�e�d�d�f�l�F��H����V��^�E��w�u�u�u�d�l�W���[����W��_�D��e�e�e�e�g�m�G��[��ƹF� \�H���e�d�d�d�g�l�F��I����W��^�D��y�_�u�u�`�l�J���I����W��_�D��d�d�e�d�f�l�G��U���F��\��K���e�d�d�d�f�l�F��H����W��_�D���u�u�u�f�e�}�I���I����W��_�E��d�e�d�d�f�l�G���Y���U��N��U��d�d�d�e�f�l�G��H����V��_�D���_�u�u�b�b�`�W��H����V��_�D��e�e�d�d�g�l�G��s��� Q��S�W��d�d�d�d�f�l�F��I����W��_�W���u�u�f�g�w�c�U��H����W��_�E��e�e�d�d�f�l�U���Y���T��
P��E��d�d�e�d�f�m�G��I����W��^�Y�ߊu�u�b�l�j�}�G��H����W��^�D��d�d�d�d�f�m�[�ԜY���� V�	N��E��d�d�d�d�f�l�F��I����V��^��U���u�f�f�u�i��G��H����W��_�D��d�e�e�e�g��W���Y����F�L�D��d�e�d�d�g�l�G��H����V��L����u�b�f�h�w�m�F��H����W��_�E��e�e�e�e�f�q�}���Y����[�^�D��d�d�d�d�f�m�G��H����W��B��U���f�f�u�k�u�m�F��H����W��^�D��d�d�d�e�u�}�W���J����X�^�D��e�d�d�e�f�m�G��I����W��NךU���b�b�h�u�g�l�F��I����V��^�E��d�e�e�e�{�W�W���N���F�_�D��d�d�d�d�g�l�F��H����V�d��U��f�u�k�w�g�l�F��H����W��_�D��e�e�e�w�w�}�W��M���D��_�D��d�d�e�d�g�l�F��H����D�=N��U��d�h�u�e�f�l�F��H����W��^�D��d�e�d�y�]�}�W��K���V��_�D��d�d�d�e�g�l�F��I����J�N��F��u�k�w�e�f�l�F��H����V��^�E��d�e�w�u�w�}�D��Y���V��_�E��d�e�d�d�f�l�F��H����FǻN��B���h�u�e�d�f�l�G��H����W��_�E��d�e�y�_�w�}�@��D���W��_�D��d�d�e�d�g�m�G��I���l�N�A���k�w�e�d�f�l�F��H����W��_�D��d�w�u�u�w�n�C���G����W��_�D��e�d�d�d�g�m�G��I���9F�]�L��u�e�d�d�f�m�F��I����W��_�D��e�y�_�u�w�j�G��Y����W��^�D��d�e�d�d�f�l�G��H���F�Y�U��w�e�d�d�f�l�F��H����V��^�D��w�u�u�u�d�h�W���[����W��_�D��d�e�e�d�f�m�F��[��ƹF� [�H���e�d�d�d�g�l�F��H����V��^�E��y�_�u�u�`�i�J���I����W��_�D��d�e�d�d�g�m�F��U���F��[��K���e�d�d�d�f�l�F��H����V��^�E���u�u�u�f�b�}�I���I����W��_�E��e�e�d�d�f�m�F���Y���U�� N��U��d�d�d�e�f�l�G��I����W��^�D���_�u�u�b�o�`�W��H����V��_�D��d�e�e�e�f�l�G��s��� Q��S�W��d�d�d�d�f�l�F��H����W��_�W���u�u�f�c�w�c�U��H����W��_�D��e�e�d�d�g�m�U���Y���P��
P��E��d�d�e�d�f�m�F��I����W��_�Y�ߊu�u�b�g�j�}�G��H����W��^�D��d�d�e�e�g�l�[�ԜY����U�	N��E��d�d�d�d�f�l�F��I����W��^��U���u�f�c�u�i��G��H����W��_�D��e�d�e�d�g��W���Y����F�L�D��d�e�d�d�g�l�F��I����W��L����u�b�c�h�w�m�F��H����W��_�D��d�d�e�d�f�q�}���Y����[�^�D��d�d�d�d�f�l�F��H����V��B��U���f�c�u�k�u�m�F��H����W��_�D��e�d�d�e�u�}�W���J����X�^�D��e�d�d�e�f�l�F��I����W��NךU���b�e�h�u�g�l�F��I����W��^�E��e�e�e�e�{�W�W���N���F�_�D��d�d�d�e�g�m�G��I����W�d��U��b�u�k�w�g�l�F��H����V��^�D��e�e�d�w�w�}�W��N���D��_�D��d�d�d�e�g�l�G��I����D�=N��U��a�h�u�e�f�l�F��H����V��_�E��d�d�d�y�]�}�W��L���V��_�D��d�d�e�e�f�m�G��I����J�N��F��u�k�w�e�f�l�F��H����V��^�E��e�e�w�u�w�}�D��Y���V��_�E��d�d�e�e�g�l�G��I����FǻN��B��h�u�e�d�f�l�G��H����V��^�D��d�e�y�_�w�}�@��D���W��_�D��d�e�e�d�f�m�F��I���l�N�M���k�w�e�d�f�l�F��H����W��_�E��d�w�u�u�w�n�O���G����W��_�D��d�e�d�e�f�m�F��H���9F�]�G��u�e�d�d�f�m�F��H����V��^�E��d�y�_�u�w�j�D��Y����W��^�D��e�e�e�e�g�l�F��H���F�Y�U��w�e�d�d�f�l�F��I����V��_�E��w�u�u�u�d�e�W���[����W��_�D��e�d�d�d�g�l�G��[��ƹF� V�H���e�d�d�d�g�l�F��I����V��_�D��y�_�u�u�`�j�J���I����W��_�D��e�d�d�e�f�m�F��U���F��V��K���e�d�d�d�f�l�F��I����W��_�D���u�u�u�f�o�}�I���I����W��_�D��d�d�d�e�g�m�F���Y���U��N��U��d�d�d�e�f�l�F��H����V��^�E���_�u�u�b�f�`�W��H����V��_�E��e�e�e�e�f�l�G��s��� Q��S�W��d�d�d�d�f�l�G��I����V��^�W���u�u�f�l�w�c�U��H����W��_�E��e�d�e�e�f�l�U���Y���_��
P��E��d�d�e�d�f�l�G��H����W��_�Y�ߊu�u�b�`�j�}�G��H����W��_�D��e�d�d�d�f�m�[�ԜY����
P�	N��E��d�d�d�d�f�m�F��H����V��_��U���u�f�l�u�i��G��H����W��^�E��e�d�d�e�f��W���Y����F�L�D��d�e�d�d�f�m�G��I����V��L����u�b�l�h�w�m�F��H����W��^�D��d�d�d�d�g�q�}���Y����[�^�D��d�d�d�d�g�l�F��I����V��B��U���f�e�u�k�u�m�F��H����W��_�D��e�e�e�e�u�}�W���J����X�^�D��e�d�d�d�g�m�F��H����V��NךU���m�f�h�u�g�l�F��I����W��_�E��e�d�d�d�{�W�W���A���F�_�D��d�d�d�e�f�m�F��I����V�d��U��e�u�k�w�g�l�F��H����V��^�E��e�e�e�w�w�}�W��I���D��_�D��d�d�d�e�f�l�F��H����D�=N��U��b�h�u�e�f�l�F��H����V��_�D��e�e�e�y�]�}�W��A���V��_�D��d�d�e�d�f�m�G��H����J�N��F��u�k�w�e�f�l�F��H����W��^�E��e�e�w�u�w�}�D��Y���V��_�E��d�d�e�d�g�l�G��I����FǻN��M��h�u�e�d�f�l�G��H����W��^�D��d�e�y�_�w�}�O��D���W��_�D��d�e�d�d�g�l�G��I���l�N�D���k�w�e�d�f�l�F��H����W��^�D��d�w�u�u�w�n�F���G����W��_�D��d�d�e�e�g�m�F��H���9F�]�@��u�e�d�d�f�m�F��H����V��_�D��e�y�_�u�w�e�A��Y����W��^�D��e�e�e�d�g�m�G��H���F�V�U��w�e�d�d�f�l�F��I����V��^�D��w�u�u�u�d�l�W���[����W��_�D��d�e�d�d�f�l�F��[��ƹF�_�H���e�d�d�d�g�l�F��H����W��^�D��y�_�u�u�o�m�J���I����W��_�D��e�d�e�d�g�l�F��U���F��_��K���e�d�d�d�f�l�F��I����W��^�E���u�u�u�f�e�}�I���I����W��_�D��e�e�d�d�g�l�G���Y���U��N��U��d�d�d�e�f�l�F��I����V��_�D���_�u�u�m�c�`�W��H����V��_�E��d�e�d�d�g�m�F��s��� ^��S�W��d�d�d�d�f�l�G��H����W��_�W���u�u�f�g�w�c�U��H����W��_�D��e�e�e�e�g�m�U���Y���T��
P��E��d�d�e�d�f�l�F��I����V��_�Y�ߊu�u�m�m�j�}�G��H����W��_�E��d�e�e�e�f�l�[�ԜY����_�	N��E��d�d�d�d�f�m�G��I����V��^��U���u�f�f�u�i��G��H����W��^�D��d�e�e�e�g��W���Y����F�L�D��d�e�d�d�f�l�F��I����W��L����u�m�g�h�w�m�F��H����W��_�D��e�d�e�e�f�q�}���Y����[�^�D��d�d�d�d�g�m�F��I����V��B��U���f�f�u�k�u�m�F��H����W��^�E��e�d�d�e�u�}�W���J����X�^�D��e�d�d�d�f�l�G��H����V��NךU���m�c�h�u�g�l�F��I����W��_�E��d�d�d�d�{�W�W���A���F�_�D��d�d�d�e�g�l�F��H����V�d��U��f�u�k�w�g�l�F��H����V��_�D��d�d�d�w�w�}�W��J���D��_�D��d�d�d�d�g�m�G��H����D�=N��U��e�h�u�e�f�l�F��H����W��^�E��e�d�d�y�]�}�W��H���V��_�D��d�d�e�d�g�l�G��I����J�N��F��u�k�w�e�f�l�F��H����W��^�E��e�e�w�u�w�}�D��Y���V��_�E��d�d�d�e�f�l�F��I����FǻN��M��h�u�e�d�f�l�G��H����V��_�E��d�e�y�_�w�}�O��D���W��_�D��d�e�d�d�g�m�G��I���l�N�A���k�w�e�d�f�l�F��H����W��_�E��e�w�u�u�w�n�C���G����W��_�D��d�d�e�e�g�m�F��H���9F�]�M��u�e�d�d�f�m�F��H����V��_�D��e�y�_�u�w�e�N��Y����W��^�D��e�d�d�e�g�m�F��H���F�V�U��w�e�d�d�f�l�F��I����W��^�E��w�u�u�u�d�h�W���[����W��_�D��d�e�d�d�f�l�G��[��ƹF�[�H���e�d�d�d�g�l�F��H����V��^�D��y�_�u�u�o�n�J���I����W��_�D��d�e�e�d�g�m�F��U���F��Z��K���e�d�d�d�f�l�F��H����W��_�E���u�u�u�f�b�}�I���I����W��_�D��d�d�e�e�g�l�G���Y���U��N��U��d�d�d�e�f�l�F��H����W��_�D���_�u�u�m�`�`�W��H����V��_�E��e�d�e�d�g�m�F��s��� ^��S�W��d�d�d�d�f�l�G��I����V��_�W���u�u�f�`�w�c�U��H����W��_�D��e�e�d�e�g�m�U���Y���P��
P��E��d�d�e�d�f�l�F��I����V��_�Y�ߊu�u�m�d�j�}�G��H����W��_�D��d�e�e�e�g�l�[�ԜY����T�	N��E��d�d�d�d�f�m�F��I����V��_��U���u�f�c�u�i��G��H����W��^�D��d�d�e�d�g��W���Y����F�L�D��d�e�d�d�f�l�F��I����W��L����u�m�`�h�w�m�F��H����W��_�D��d�e�e�d�g�q�}���Y����[�^�D��d�d�d�d�f�m�G��H����W��B��U���f�c�u�k�u�m�F��H����W��^�E��e�d�e�e�u�}�W���J����X�^�D��e�d�d�d�g�m�G��H����V��NךU���m�l�h�u�g�l�F��I����W��^�D��d�d�d�d�{�W�W���A���F�_�D��d�d�d�d�g�m�G��I����W�d��U��b�u�k�w�g�l�F��H����W��^�E��d�d�d�w�w�}�W��N���D��_�D��d�d�d�e�g�l�F��I����D�=N��U��f�h�u�e�f�l�F��H����V��^�E��d�d�d�y�]�}�W��M���V��_�D��d�d�d�e�f�m�G��I����J�N��F��u�k�w�e�f�l�F��H����V��_�D��e�e�w�u�w�}�D��Y���V��_�E��d�d�e�e�g�l�F��I����FǻN��M��h�u�e�d�f�l�G��H����V��^�E��e�d�y�_�w�}�O��D���W��_�D��d�d�e�d�g�l�G��H���l�N�B���k�w�e�d�f�l�F��H����W��_�D��e�w�u�u�w�n�O���G����W��_�D��d�e�e�d�f�m�G��I���9F�]�D��u�e�d�d�f�m�F��H����V��^�D��e�y�_�u�w�e�E��Y����W��^�D��d�e�e�e�f�l�G��H���F�V�U��w�e�d�d�f�l�F��H����W��_�D��w�u�u�u�d�e�W���[����W��_�D��e�d�e�d�f�m�G��[��ƹF�V�H���e�d�d�d�g�l�F��I����V��^�E��y�_�u�u�o�k�J���I����W��_�D��e�e�e�d�g�l�F��U���F��Y��K���e�d�d�d�f�l�F��I����W��_�E���u�u�u�f�o�}�I���I����W��_�D��d�d�d�d�g�l�G���Y���U��N��U��d�d�d�e�f�l�F��H����W��_�D���_�u�u�m�g�`�W��H����V��_�D��d�e�d�e�f�m�G��s��� ^��S�W��d�d�d�d�f�l�F��H����V��_�W���u�u�f�l�w�c�U��H����W��_�E��e�d�d�e�f�m�U���Y���_��
P��E��d�d�e�d�f�l�G��H����V��_�Y�ߊu�u�m�a�j�}�G��H����W��_�E��e�d�d�d�f�l�[�ԜY����
S�	N��E��d�d�d�d�f�l�G��H����V��^��U���u�f�l�u�i��G��H����W��_�D��d�e�e�e�g��W���Y����F�L�D��d�e�d�d�f�m�G��I����V��L����u�m�m�h�w�m�F��H����W��^�E��d�e�e�e�f�q�}���Y����[�^�D��d�d�d�d�f�l�G��H����V��B��U���f�e�u�k�u�m�F��H����W��_�E��d�d�e�e�u�}�W���J����X�^�D��e�d�d�d�g�m�F��H����W��NךU���l�g�h�u�g�l�F��I����W��^�E��e�d�d�e�{�W�W���@���F�_�D��d�d�d�d�f�m�F��I����W�d��U��e�u�k�w�g�l�F��H����W��^�D��d�d�e�w�w�}�W��I���D��_�D��d�d�d�e�g�m�G��I����D�=N��U��c�h�u�e�f�l�F��H����V��^�E��d�e�d�y�]�}�W��N���V��_�D��d�d�d�d�f�m�F��I����J�N��F��u�k�w�e�f�l�F��H����W��_�D��d�d�w�u�w�}�D��Y���V��_�E��d�d�e�e�g�l�F��H����FǻN��L��h�u�e�d�f�l�G��H����V��^�D��e�d�y�_�w�}�N��D���W��_�D��d�d�d�d�g�l�G��I���l�N�D���k�w�e�d�f�l�F��H����W��^�D��e�w�u�u�w�n�F���G����W��_�D��d�e�e�d�f�l�F��H���9F�]�A��u�e�d�d�f�m�F��H����V��^�E��d�y�_�u�w�d�B��Y����W��^�D��d�d�e�e�g�m�G��H���F�W�U��w�e�d�d�f�l�F��H����V��_�D��w�u�u�u�d�l�W���[����W��_�D��e�d�e�e�f�l�G��[��ƹF�_�H���e�d�d�d�g�l�F��I����W��^�D��y�_�u�u�n�d�J���I����W��_�D��d�e�e�d�g�l�F��U���F��^��K���e�d�d�d�f�l�F��H����V��^�D���u�u�u�f�e�}�I���I����W��_�D��d�d�e�e�f�l�G���Y���U��N��U��d�d�d�e�f�l�F��H����V��^�E���_�u�u�l�d�`�W��H����V��_�D��e�d�d�d�f�m�G��s��� _��S�W��d�d�d�d�f�l�F��H����W��^�W���u�u�f�g�w�c�U��H����W��_�E��e�d�e�d�g�l�U���Y���
T��
P��E��d�d�e�d�f�l�G��I����V��_�Y�ߊu�u�l�b�j�}�G��H����W��_�D��d�e�d�e�g�l�[�ԜY����^�	N��E��d�d�d�d�f�l�F��I����V��^��U���u�f�g�u�i��G��H����W��_�D��e�d�d�e�g��W���Y����F�L�D��d�e�d�d�f�m�F��H����V��L����u�l�d�h�w�m�F��H����W��^�D��e�d�d�e�g�q�}���Y����[�^�D��d�d�d�d�f�l�F��I����W��B��U���f�f�u�k�u�m�F��H����W��^�E��e�e�e�e�u�}�W���J����X�^�D��e�d�d�d�f�m�G��H����V��NךU���l�`�h�u�g�l�F��I����W��^�E��e�d�d�d�{�W�W���@���F�_�D��d�d�d�d�g�m�F��I����W�d��U��f�u�k�w�g�l�F��H����W��^�D��d�e�e�w�w�}�W��J���D��_�D��d�d�d�d�g�m�F��H����D�=N��U��l�h�u�e�f�l�F��H����W��_�D��e�e�e�y�]�}�W��I���V��_�D��d�d�d�e�g�m�G��I����J�N��F��u�k�w�e�f�l�F��H����V��_�E��e�e�w�u�w�}�D��Y���V��_�E��d�d�d�e�f�m�F��H����FǻN��L��h�u�e�d�f�l�G��H����V��_�E��e�d�y�_�w�}�N��D���W��_�D��d�d�e�d�g�m�G��I���l�N�A���k�w�e�d�f�l�F��H����W��^�D��d�w�u�u�w�n�C���G����W��_�D��d�d�e�e�f�l�G��I���9F�]�B��u�e�d�d�f�m�F��H����V��^�E��e�y�_�u�w�d�O��Y����W��^�D��d�e�d�d�g�l�F��I���F�W�U��w�e�d�d�f�l�F��H����W��_�E��w�u�u�u�d�h�W���[����W��_�D��d�e�d�e�g�m�F��[��ƹF�[�H���e�d�d�d�g�l�F��H����W��_�D��y�_�u�u�n�o�J���I����W��_�D��e�d�d�e�g�l�G��U���F��]��K���e�d�d�d�f�l�F��I����W��_�D���u�u�u�f�b�}�I���I����W��_�D��e�d�d�d�g�l�F���Y���U��N��U��d�d�d�e�f�l�F��H����V��^�D���_�u�u�l�a�`�W��H����V��_�D��e�e�d�e�f�m�F��s��� _��S�W��d�d�d�d�f�l�F��I����W��^�W���u�u�f�`�w�c�U��H����W��_�D��e�e�e�d�f�l�U���Y���
S��
P��E��d�d�e�d�f�l�F��I����V��_�Y�ߊu�u�l�e�j�}�G��H����W��_�E��d�e�d�e�g�l�[�ԜY����W�	N��E��d�d�d�d�f�l�G��I����W��_��U���u�f�c�u�i��G��H����W��_�D��e�e�d�d�g��W���Y���� F�L�D��d�e�d�d�f�l�F��H����V��L����u�l�a�h�w�m�F��H����W��_�E��e�e�e�d�f�q�}���Y����[�^�D��d�d�d�d�f�m�G��H����V��B��U���f�c�u�k�u�m�F��H����W��^�D��d�e�e�d�u�}�W���J����X�^�D��e�d�d�d�f�l�F��H����W��NךU���l�m�h�u�g�l�F��I����W��_�E��e�e�d�d�{�W�W���@���F�_�D��d�d�d�d�g�l�G��H����V�d��U��b�u�k�w�g�l�F��H����W��_�D��e�e�d�w�w�}�W��N���D��_�D��d�d�d�d�f�m�G��H����D�=N��U��g�h�u�e�f�l�F��H����W��^�D��e�e�e�y�]�}�W��J���V��_�D��d�d�d�e�f�l�F��H����J�N��F��u�k�w�e�f�l�F��H����V��^�E��d�e�w�u�w�}�D��Y���V��_�E��d�d�d�d�f�m�G��I����FǻN��L��h�u�e�d�f�l�G��H����W��_�E��d�e�y�_�w�}�N��D���W��_�D��d�d�e�d�g�l�F��H���l�N�B���k�w�e�d�f�l�F��H����W��^�D��e�w�u�u�w�n�@���G����W��_�D��d�d�d�d�f�m�G��H���9F�]�E��u�e�d�d�f�m�F��H����W��^�E��e�y�_�u�w�d�F��Y����W��^�D��d�d�e�e�g�l�G��H���F�W�U��w�e�d�d�f�l�F��H����V��_�E��w�u�u�u�d�e�W���[����W��_�D��d�e�e�d�g�l�F��[��ƹF�V�H���e�d�d�d�g�l�F��H����W��^�D��y�_�u�u�n�h�J���I����W��_�D��d�e�d�e�g�m�G��U���F��X��K���e�d�d�d�f�l�F��H����W��_�D���u�u�u�f�o�}�I���I����W��_�D��e�e�d�d�g�m�G���Y���U��N��U��d�d�d�e�f�l�F��I����W��_�E���_�u�u�l�n�`�W��H����V��_�D��e�e�e�d�f�l�F��s��� _��S�W��d�d�d�d�f�l�F��I����W��_�W���u�u�f�l�w�c�U��H����W��_�D��d�d�d�d�g�m�U���Y���
_��
P��E��d�d�e�d�f�l�F��H����W��_�Y�ߊu�u�l�f�j�}�G��H����W��_�D��d�e�d�e�g�l�[�ԜY����
R�	N��E��d�d�d�d�f�l�F��H����W��^��U���u�f�l�u�i��G��H����W��_�E��d�d�e�d�g��W���Y����F�L�D��d�e�d�d�f�l�G��H����V��L����u�l�b�h�w�m�F��H����W��_�D��e�d�e�d�g�q�}���Y����[�^�D��d�d�d�d�f�l�F��H����V��B��U���f�l�u�k�u�m�F��H����W��_�E��d�d�d�e�u�}�W���M����X�^�D��e�d�d�d�f�m�G��H����W��NךU���e�d�h�u�g�l�F��I����W��^�D��e�e�e�d�{�W�W���I���F�_�D��d�d�d�d�f�l�F��H����V�d��U��e�u�k�w�g�l�F��H����W��_�D��e�e�d�w�w�}�W��I���D��_�D��d�d�d�d�g�m�F��H����D�=N��U��`�h�u�e�f�l�F��H����W��_�E��d�e�d�y�]�}�W��O���V��_�D��d�d�d�d�f�m�G��H����J�N��A��u�k�w�e�f�l�F��H����W��^�D��e�e�w�u�w�}�C��Y���V��_�E��d�d�d�e�f�l�F��H����FǻN��E��h�u�e�d�f�l�G��H����V��_�E��d�d�y�_�w�}�G��D���W��_�D��d�d�d�d�f�m�F��H���l�N�D���k�w�e�d�f�l�F��H����W��_�D��d�w�u�u�w�i�F���G����W��_�D��d�d�e�d�f�m�G��I���9F�Z�F��u�e�d�d�f�m�F��H����W��_�E��e�y�_�u�w�m�C��Y����W��^�D��d�d�d�d�f�m�F��H���F�^�U��w�e�d�d�f�l�F��H����V��_�E��w�u�u�u�c�l�W���[����W��_�D��d�d�e�e�g�l�F��[��ƹF�_�H���e�d�d�d�g�l�F��H����V��_�D��y�_�u�u�g�e�J���I����W��_�D��d�e�e�e�g�m�F��U���F��W��K���e�d�d�d�f�l�F��H����W��^�D���u�u�u�a�e�}�I���I����W��_�D��d�e�e�e�f�l�F���Y���R��N��U��d�d�d�e�f�l�F��H����W��^�D���_�u�u�e�e�`�W��H����V��_�D��e�d�d�e�f�l�F��s���V��S�W��d�d�d�d�f�l�F��I����W��^�W���u�u�a�g�w�c�U��H����W��_�D��e�d�e�e�g�m�U���Y���T��
P��E��d�d�e�d�f�l�F��I����W��^�Y�ߊu�u�e�c�j�}�G��H����W��_�D��e�e�d�e�g�l�[�ԜY����Q�	N��E��d�d�d�d�f�l�F��I����V��_��U���u�a�g�u�i��G��H����W��_�D��e�d�d�d�g��W���Y����
F�L�D��d�e�d�d�f�l�F��H����W��L����u�e�e�h�w�m�F��H����W��_�E��d�e�e�e�g�q�}���Y����[�^�D��d�d�d�d�f�l�G��H����W��B��U���a�f�u�k�u�m�F��H����W��_�D��e�e�e�d�u�}�W���M����X�^�D��e�d�d�d�f�l�F��H����V��NךU���e�a�h�u�g�l�F��I����W��_�D��d�d�e�e�{�W�W���I���F�_�D��d�d�d�d�f�m�F��I����V�d��U��f�u�k�w�g�l�F��H����W��^�D��d�e�d�w�w�}�W��J���D��_�D��d�d�d�d�f�l�F��H����D�=N��U��m�h�u�e�f�l�F��H����W��_�D��e�e�e�y�]�}�W��@���V��_�D��d�d�d�d�f�m�G��H����J�N��A��u�k�w�e�f�l�F��H����W��^�D��e�d�w�u�w�}�C��Y���V��_�E��d�d�d�d�g�m�G��H����FǻN��E��h�u�e�d�f�l�G��H����W��^�D��e�d�y�_�w�}�G��D���W��_�D��d�d�d�d�g�m�F��H���l�N�A���k�w�e�d�f�l�F��H����W��^�D��e�w�u�u�w�i�C���G����W��_�D��d�d�d�e�f�m�F��H���9F�Z�C��u�e�d�d�f�m�F��H����V��_�D��e�y�_�u�w�m�@��Y����W��^�D��d�d�d�d�g�l�G��I���F�^�U��w�e�d�d�f�l�F��H����W��_�E��w�u�u�u�c�i�W���[����W��_�D��d�d�e�e�g�m�F��[��ƹF�[�H���e�d�d�d�g�l�F��H����V��^�D��y�_�u�u�g�l�J���I����W��_�D��d�d�d�e�g�l�F��U���F��\��K���e�d�d�d�f�l�F��H����V��^�E���u�u�u�a�b�}�I���I����W��_�D��d�e�d�e�g�m�F���Y���R��N��U��d�d�d�e�f�l�F��H����W��^�E���_�u�u�e�b�`�W��H����V��_�D��d�d�d�d�g�l�G��s���V��S�W��d�d�d�d�f�l�F��H����W��^�W���u�u�a�`�w�c�U��H����W��_�D��d�e�d�d�f�m�U���Y���S��
P��E��d�d�e�d�f�l�F��H����V��_�Y�ߊu�u�e�l�j�}�G��H����W��_�D��e�d�d�e�f�l�[�ԜY����V�	N��E��d�d�d�d�f�l�F��I����V��_��U���u�a�c�u�i��G��H����W��_�D��d�e�e�d�g��W���Y����F�L�D��d�e�d�d�f�l�F��H����W��L����u�e�f�h�w�m�F��H����W��_�D��e�d�e�e�f�q�}���Y����[�^�D��d�d�d�d�f�l�F��H����V��B��U���a�c�u�k�u�m�F��H����W��_�D��e�e�d�d�u�}�W���M����X�^�D��e�d�d�d�f�l�F��H����W��NךU���e�b�h�u�g�l�F��I����W��_�E��d�d�e�e�{�W�W���I���F�_�D��d�d�d�d�f�l�F��I����W�d��U��c�u�k�w�g�l�F��H����W��_�E��d�d�e�w�w�}�W��N���D��_�D��d�d�d�d�f�l�G��H����D�=N��U��d�h�u�e�f�l�F��H����W��_�E��d�d�d�y�]�}�W��K���V��_�D��d�d�d�d�f�l�F��H����J�N��A��u�k�w�e�f�l�F��H����W��_�E��e�d�w�u�w�}�C��Y���V��_�E��d�d�d�d�f�m�F��H����FǻN��E���h�u�e�d�f�l�G��H����W��^�D��e�e�y�_�w�}�G��D���W��_�D��d�d�d�d�f�m�G��I���l�N�B���k�w�e�d�f�l�F��H����W��^�E��d�w�u�u�w�i�@���G����W��_�D��d�d�d�d�f�m�F��I���9F�Z�L��u�e�d�d�f�m�F��H����W��_�D��d�y�_�u�w�m�G��Y����W��^�D��d�d�d�d�g�l�G��I���F�^�U��w�e�d�d�f�l�F��H����W��_�D��w�u�u�u�c�e�W���[����W��_�D��d�d�d�d�g�m�F��[��ƹF�V�H���e�d�d�d�g�l�F��H����W��_�E��y�_�u�u�g�i�J���I����W��_�D��d�d�d�d�f�m�F��U���F��[��K���e�d�d�d�f�l�F��H����W��^�D���u�u�u�a�o�}�I���I����W��_�D��d�d�d�d�g�m�G���Y���R�� N��U��d�d�d�e�f�l�F��H����W��_�E���_�u�u�e�o�`�W��H����V��_�D��d�d�d�e�f�m�F��s���V��S�W��d�d�d�d�f�l�F��H����W��_�W���u�u�a�l�w�c�U��H����W��_�D��d�d�d�e�g�m�U���Y���_��
P��E��d�d�e�d�f�l�F��H����W��^�Y�ߊu�u�e�g�j�}�G��H����W��_�D��d�d�d�e�f�m�[�ԜY����
U�	N��E��d�d�d�d�f�l�F��H����W��_��U���u�a�l�u�i��G��H����W��_�D��d�d�d�d�f��W���Y����F�L�D��d�e�d�d�f�l�F��H����W��L����u�e�c�h�w�m�F��H����V��^�E��e�e�e�e�g�}�L�Զ����Q��+��<���������(���6����	F��E��N��2�;�_�_�2�2��������T��S1�U���6�&�u�4�3�m�W����ƹF���ڊ�8�u�h�4�3�m�}��� ����@��C�����0�:�3�u�w�}����:����z(��p+�����e�u�u�0��4���Y����9F�N��U���4�1�e�!�'�a�WǱ�����X�I����u�u�9�0�]�}�W���Y����W��h��U��4�1�e�_�w�}�W���Y����K��Y�����!�4�&�4�2�2�}���Y����V��=d�����4�6�&�o�'�2����Q����F��R	��U���u�<�u�6�<�8��������_�I�\ʡ�0�_�u�u�w�}�������W����ߊu�u�u�u�w�}�G��Y����p)��h'��0���}�1�'�
�:�t�L�ԜY���F��SN��N���u�0�1�<�l�8�Ϯ�����l��Y
����_��7�4�.��2������v#��D�����6�d�c�{�;�f�}�������uR��/����3�l�>�'��}����YӁ��V��FךU���u�u�4�4�>�)�W���7����aF��]����u�u�u�1�%�.�%�������}2��r<��H��l�n�u�u�w�}�6�������W��N��!����o�u�f�l�}�WϮ����F�N�����!�o��u���8���B���F���U���������}���Y���R��R��U���������!���6�΍�W��D9�����u�u����m�L���Y�����T��;ʆ�����]�}�W���Y���)��=��*����
�����������W��x9��:��|�_�;�u�9�4��Զ����G��B�����u�3�8�a�a��O���&����X��hX�����u�6�8�:�2�)���Oʧ��U9��Q1�����
�
�:�u�$�}�W���YӖ��GF�N��U���u�u�6�>�m��W���&����p]ǻN��U���u�u�1�'�w�}�9ύ�=����z%��r-��'�ߊu�u�u�u�w�}����Y����g"��x)��N���u�u�u�u�w�,�W���,�Ɵ�w9��p'��#����|�_�u�w�3�W���	����G]Ǒ=d�����u�u�8�a�a��O���&����X��hX�����u�u�6�8�8�8�ϳ�M���� ^��1��L���'�
�
�:�]�}�W���Ӌ��NǻN��U���9�u�k�6�<�W�W���Y�ƭ�W��
P�����&�e�_�u�w�}�W���Y����VV�N��U���$�u�k�$�~�W��������G��B����