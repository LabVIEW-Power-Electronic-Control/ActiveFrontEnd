-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�a�c��m���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����V��Y1�Oʚ�������!���6���F��@ ��U���_�u�u�%�%�)����Y�ƃ�gF��s1��2������u�d�}�������9F������u������4���s����9l��E����� �0�7�=�!�2�W���I�ߍ� ��h��U���_�u�u�:�$�<�Ͽ�&����G9��P��D�������g�W��B�����D��ʴ�
�:�&�
�8�4�(���Y����)��tN�U��n�u�u�6�9�)����	����@��Q��E��������4���Y����\��XN�U��w�e�d�n�w�}��������R��c1��G���8�d�o����0���/����aF�
�����e�u�h�w�g�m�L���YӅ��@��CN��*���&�f�3�8�e�g�$���5����l0��c!��]���:�;�:�e�w�`�U��I��ƹF��X �����4�
��&�c�;���Cӵ��l*��~-��0����}�u�:�9�2�G���D����V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����F��d:��9�������w�m��������\�_�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��d�w�_�u�w�2����Ӈ��P	��C1��F؊��o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�d�d�n�w�}��������R��X ��*���g�f�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�d�e�e�u�W�W�������]��G1�����9�f�
��m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�d�f�m�L���YӅ��@��CN��*���&�
�#�a�g�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��Cي�u�u��
���(���-���T��X����u�h�w�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��D؊�f�u�u����>���<����N��
�����e�u�h�w�f�m�G��I���9F������!�4�
�:�$�����=����g"��x)��*�����}�d�3�*����P���V��^�E��d�n�u�u�4�3����Y����\��h��G���f�o�����4���:����W��S�����|�o�u�d�f�l�F��H����F�T�����u�%�6�;�#�1�F݁�O����g"��x)��*�����}�d�3�*����P���V��^�D��e�n�u�u�4�3����Y����\��h��G���o������!���6���F��@ ��U���o�u�e�e�g�m�F��[���F��Y�����%�6�;�!�;�l�(ܘ�?����g"��x)��*�����}�f�3�*����P���W��_�D��d�d�n�u�w�>�����ƭ�l��D�����e�o�����4���:����W��S�����|�o�u�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����	F��s1��2������u�f�}�������	[�_�D��e�d�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�e�w�]�}�W���
������T�����d�
�e�d�m��3���>����v%��eN��Fʱ�"�!�u�|�m�}�G��I����V��L�U���6�;�!�;�w�-�������� 9��N��1��������}�F�������V�S��E��e�e�e�e�g�f�W�������R��V�����
�#�f�d�g�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�N���u�6�;�!�9�}��������EW��^�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��G��I���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=d��Uʦ�2�4�u�%������Y����)��t1��6���u�f�1�"�#�}�^��Y����D��N�����<� �0�3�:�8��������@��Y	�U���4�!�<� �2�;��������TF����6���&�u�u�<�9�1��������l�N�����u�%�&�2�4�8�(���
�ד�@��T��!�����n�u�w�.����Y����Z��S
��G������]�}�W�������R��1�����&�u�u����>���<����N��
�����e�n�u�u�$�:��������l��T��!�����n�u�w�.����Y����lP��N�&���������W��Y����G	�UךU���<�;�9�%��1�(ځ�����l��N��1��������}�F�������V�=N��U���;�9�%��;��(���&����	F��s1��2������u�f�}�������9F������!�%�g�
�2��E���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T���������!�g��(�C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���9�-���#�o�(���&����	F��s1��2������u�g�9� ���Y����F�D�����%�&�2�6�2��#���K����lW�=��*����n�u�u�$�:����	����l��h[�Oʗ����_�w�}����ӓ��K5��N!��*���3�
�a�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������O=�����
�f�'�2�b�d�Mύ�=����z%��r-��'���g�1�"�!�w�t�}���Y����R
��d1��1����!�'�
�o�4��������R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�3���2���+����lU��^ �����'�2�`�`�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƪ�l/��r6��'���8�a�
�;�6�:�(���M�ߓ�F��d:��9�������w�m��������l�N�����u���������&�ד�]��P�����`�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�&����P��h=�����3�8�g�o���;���:���F��P ��U���&�2�7�1�`�}�W���5����9F������3�
����(�(�������F��d:��9�������w�n�W������]ǻN�����9�3�
���	����H����l ��^�����u��
����2���+������Y��E��u�u�&�2�6�}�$���5����F��1����d�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�&����P��h=�����3�8�f�o���;���:���F��P ��U���&�2�7�1�n�}�W���5����9F������!�%�d�
�"�i�C���Y�Ɵ�w9��p'��#����u�c�u�8�3���B�����Y�����d�
� �a�c�-�W���-����t/��a+��:���c�u�:�;�8�m�L���Yӕ��]��S1�����
� �d�f�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��R	��*���d�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ʃ�C9��G1�����f�
�a�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lW��Q��A݊�d�o�����4���:����S��S�����|�_�u�u�>�3�Ϫ�	����S��G]��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u��8����
����S��G_��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�$�8�(���H�ӓ� F��d:��9�������w�m��������l�N�����u�4�
�
��(�F���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʡ�%�b�3�
�e��F��*����|!��h8��!���}�g�1�"�#�}�^�ԜY�ƿ�T����*ӊ� �d�f�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����uT��B1�F���u�u��
���(���-���W��X����n�u�u�&�0�<�W���&����lW��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��(���H�ӓ�F��d:��9�������w�l�W������]ǻN�����9�!�%�`�1��Gށ�K����g"��x)��*�����}�d�3�*����P���F��P ��U���4�!�3�
�g��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������g�3�
�c��n�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��_1�����&�
� �g�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��G���
�a�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������^��1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������9��h\�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����H¹��lT��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�F݁�����l��N��1��������}�D�������V�=N��U���;�9�!�%�o�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�g�
� �e�l����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N�����
�`�
�f�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������^��1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������
9��D�� ��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U��B1�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Kǹ��lU��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�5�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�d�
� �d�j����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��#���
�
� �g�`�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��C��D���
�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��Q��Dӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l ��\�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	����lU��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������T��Q��A݊�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l ��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	Ĺ��lU��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��<�E�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�0��0�D���&����CU�=��*����
����u�DϺ�����O��N�����4�u�0�
�:�l�(�������l ��Y�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)��������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-����Nʹ��\��c*��:���
�����}�������9F������&�9�!�%��(�D���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�f�3�
�`��F��*����|!��h8��!���}�f�1�"�#�}�^�ԜY�ƿ�T����*���m�3�
�c��n�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��O��0��� �
�f��1��G؁�K����g"��x)��*�����}�f�3�*����P���F��P ��U���4�g�c�3��l�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����c�3�
�g��l�Mύ�=����z%��r-��'���g�1�"�!�w�t�}���Y����R
��h8�����3�
�g�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h_�����f�
�f�o���;���:����g)��_����!�u�|�_�w�}����Ӏ��}#��x��Dӊ�:�<�!�3��k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&�����!�d��8�(���M�ԓ�F��d:��9�������w�n�W������]ǻN�����9�3�
��/�(�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u����8���Jƹ��l��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����K)��h]�����3�
�l�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��y+��:���f�
� �a�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��Q=��0���� �
�`�e�;�(��&���5��h"��<������}�f�9� ���Y����F�D����������)�Dށ�&����U��N�&���������W��Y����G	�UךU���<�;�9�4��8����I����TF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���&�2�4�u�'�/����&¹��V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�<�;�9�6��$�������g"��x)��*�����}�u�8�3���B�����Y�����<�
�1�
�g�g�5���<����F�D�����%�&�2�7�3�i�O��;����r(��N�����4�u�%�&�0�?���L����|)��v �U���&�2�4�u�'�.��������\��x!��4��_�u�u�:�'�3����?����rU��h^�����
�g�&�c��}�$���YӁ��V��FךU���u�u��o��	�0���s���F�y;��&����o�����}���Y���W��h9��!���u����l�}�W���Yӂ��G9��s:��Oʜ����|�]�}�W�����ƹF�N����o��u����>���<����N��
�����e�n�u�u�w�}����Y�ƃ�gF��s1��2������u�a�}�������]ǻN�����:�%�;�;�l�W�W�������]����E���f�3�e�3�n�6����Y��ƹF��R �����_�u�u�u�w�<��������z(��p+�����u�u�u�1�%�.�%�������}2��r<�U���u�u��1�2�.����Y�ƅ�g#��eN����u�:�!�}�w�}�W������/��d:��9����_�u�u�w�}����Y�ƅ�5��h"��<��u�u�u�u�6�9����Y�ƅ�5��h"��<������}�e�9� ���Y����F�N����o��u����>��Y���F��N�:���������4���Y����W	��C��\���_�u�u�;�w�2������Ɠ9l��P��U���>�'�
�
�w�}��������^ ��W��M���
�
�
�4�%�k�W�������Z��V�����u�u�u�4�6�4����G����9F�N��U���'�&��;�2�`�W��N���F�N�����&�<�!�u�i�l�^���YӖ��GF��GN��U���u�u�6�>�j�}�������F�N�����h�u�%�'�#�W�W���Y�ƭ�W��D^��Kʾ�'�
�
�1�%�.�G�ԜY���F��N��U���'�c�6�e�]�}�W���Y���F��E��*��n�_�u�u������&�Ԣ�lP��1��U���:�%�;�;�w��G���Jˀ��l ��O��G���c�
�_�u�w�8����Y����l�N��Uʜ�u�k�d�_�w�}�W���,����r!��
P��Y���u�u�u�1�9��>���Y���JǻN��U���:�!����`�W��s���C	����U�ߊu�u�u�u�>�m�J�������l�N��Uʱ� �u�k�1�6�.��������l��dװ�ߊu�u�x�!�2�>����ӕ��G�V��&���8�u�3�!�2�.��������]�CךU���%��
�&��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�4������E�ƭ�l(��Q�����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӇ��A��E ��*���2�4�&�2�w�/����W���F�V�����;�e�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����V��Y1�����u�h�4�
�8�.�(���K����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�!�2�}�W���Y���F�N��U���%�'�!�'������E�ƪ�l5��r-�� ���`�g�3�
�o��D�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�%�'�#�/�(ށ�����@��YN�����&�u�x�u�w�<�(�������l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�4�
�0�"�3�F��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ہ�
����O��_�����u�u�u�u�w�}�W���Y����V��Y1�����u�h�3�
���#���&�ד�l ��^����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���U5��r"��!���
�`�'�2�o�}����Ӗ��P��N����u��������&����^��D�����:�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Q����Z��S
��G���!�0�u�u�w�}�W���Y���F���&�����!�d��8�(��E�ƭ�l��D�����e�_�u�u�w�}�W���Y�Ʃ�@�������7�1�l�|�#�8�W���Y���F�N��U���u��������&����^�
N�����
�e�_�u�w�}�W���Y���V��^�U���u�u�u�u�2�9���s���F�R ����u�u�0�1�'�2����s���K�Q=��0���� �
�d�%�:�F������]F��X�����x�u�u�3���2�������l��h_�*���<�;�%�:�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y�ƥ�N��h��*���
�f�|�!�2�}�W���Y���F�N��U��������)�Dށ�����F������!�9�f�
�l�}�W���Y���F������4�
�<�
�3��G�������9F�N��U���u�u�u�u�w��$���:����lU��E��D��i�u�4�'�a�,�L���Y���F�N��U���u�3�_�u�w�}�W���Y����Z ��=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G��U���;�u�u�u�w�}�W���Yӄ��_9��r����
�0�
�f�w�`����&����|��V�� ��m�%�n�u�w�}�W���Y��� ��~ ��-���!�'�
�m�>�/��������S�
N��*������0�:�n�(�������U��V��G�ߊu�u�u�u�w�}�W���.����q��C1�*���
�f�u�h�"��$���6���� 9��hZ�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������O�C�����u�u�u�u�w�}�W���0����r4��R��Aۊ�;�4�2�
�2��B���DӀ��z(��o/�����
�d�<�'�9�8����Lʹ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�4�t�������R��C��U���%�6�;�!�;�:���P����[��N��U���u�u�u�u�'��݁�&����T��S��*���g�`�3�
�n��D�ԜY���F�N��Uʡ�%�g�
�0��o�W��	����9��Q��Lۊ�f�d�u�:�9�2�F���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p��������@��RN�����
�&�|�:�w�5�W����ơ�P��R@��X���u�4�
��1�0��������\������u�4�
�!�%�q����*����F��h�����u�0�<�_�w�}�W�������C9��h��U���u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����4�!�h�4��2��������O�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!��.�(��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�F�������F�N��U���u�u�0�1�>�f�W���Y���F��_������&�g�3�:�l�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���K����lW��N��U���u�u�u�u�2�9���Y���F�N�����4�
��&�d�;���D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&���� ]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����l ��h\�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�C������FǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�8�5����G��ƹF�N��U���u�u�%���.�W��[����]ǻN��U���;�u�4�0�]�}�W���Y����V��=N��U���3�
�m�
�e�a�W���&����P9��T��]���<�;�1�4��2�����ԓ� U�N�����0�}�8�
��(�F���	���9l�N�U���1�;�u�&�>�3�������KǻN�����;�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B�����y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Q�΢�GN��G1�����9�2�6�d�j�<�(������R�������!�9�2�6�f�`��������V��c1��D���8�e�|�:�w�u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�C������O��_�����u�u�u�u�w�-����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�:�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�3�8�����Ƽ�\��D@��X���u�4�
�1�2�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����|�u�u�7�0�3�W���Y����UF�Y��]���6�;�!�9�0�>�F������R��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�t�W������F�N��Uʴ�
�1�0�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��[��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������,�4�&�2�w�/����W���F�V�����
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&���� O����ߊu�u�u�u�w�}�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�'�4�.�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������@��YN�����&�u�x�u�w�<�(�������l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�a�3�8�d�}�$���5����F��1�����m�
�f�u�'�/����&ù��V�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���ǹ��^9��G�����_�u�u�u�w�}�W�������]9��S��&������!�f��(���M�ԓ� ]ǻN��U���9�0�_�u�w�}�W���Y����V��Y1�I���%�'�!�'������s���F�R ����_�u�u�;�w�/����B��ƹF�N��*��� �;�d�4�$�:�W�������K��N�����0� �;�d�6�.���������T��]���6�y�4�
�>�����*����9��Z1�U�������#�n�(݁�����l�������'�
�
�'�0�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^Ϫ���ƹF�N��U���%�'�!�'��}�Jϸ�&����p2��C1�*؊� �`�f�%�l�}�W���YӃ��VFǻN��U���u�u�%�'�#�/�(���DӇ��A��E ��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����W��[�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ����� ��~ ��-���!�'�
�d�>�/��������R�V�����&�$��
�#�����P�����^ ךU���u�u�u�u�w�}��������lW��R��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<�ϰ��έ�l��D��ۊ�u�u�����%�������l��V ��*���
�`�|�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(������]F��X�����x�u�u�4��4�(���&�ԓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U´�
��3�8�g�9� ���Y�����T�����d�d�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�i�OϿ�
����C��R��U���u�u�4�
�>�����K˹��@��h����%�:�0�&�6�����
����g9��1����u���������&�ޓ�]��P�� ��m�%�|�u�w�?����Y���F�N��U���%�&�2�7�3�i�O��Y�έ�l��D�����
�u�u�%�$�:����&����GT��D��\ʴ�1�}�����%�������l��V ��*���a�m�%�u�w�-��������lV�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����d�4�&�2�w�/����W���F�V�����1�
�f�
�$�4��������C��R���������2�0�Cށ�����V9��hZ�*��u�%�&�2�4�8�(���
�Փ�@��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����d�i�u�}�'�>��������lW������6�0�
��$�n����K�ƭ�WF��G1�����9�d�e�h�1��9���8����A��1�����0�3�
�`��o�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����������^	�����0�&�u�x�w�}��������W9��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��i�u�4�
�8�.�(���&���R��d1����1�"�!�u�~�f�W�������A	��D����u�x�u�%�$�:����N�ƭ�@�������{�x�_�u�w�-��������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�g�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(������]F��X�����x�u�u�4��4�(���&�֓�@��Y1�����u�'�6�&���>���!����V��V�����2�
�0�
�c�q��������V��c1��F���8�g�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��m�K���Q����\��h�����u�u�%�&�0�>����-����l ��h\�����;�!�}����/������� ^��Y�����0�
�a�u�w�-��������lV�UךU���;�u�'�6�$�f�}���Y���R��^	�����m�4�&�2�w�/����W���F�V�����1�
�m�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�d�W��Q����\��h��*���u�%��
�$�u�W������O��N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�d�3�8�g�<����Y����V��C�U���4�
�<�
�$�,�$���¹��^9��V�����'�6�o�%�8�8�ǿ�&����Q��\��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��G���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�3�8�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�f�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=�����3�8�d�4�$�:�W�������K��N�����<�
�&�$���݁�
����R��P �����o�%�:�0�$�<�(���&����P�N�����;�u�u�u�w�4�Wǿ�&����Q��X�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�d�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�g�3�:�l�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�����g�4�&�2�w�/����W���F�V�����&�$��
�#�����&����T��E��Oʥ�:�0�&�4��4�(���&���F�U�����u�u�u�<�w�<�(���&����P�C��U���u�u�u�u�w�<�(���&����l5��D�����g�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���f�3�8�g�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��Q��Fʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�
�$��(�������A	��N�����&�4�
�<��9�(��s���Q��Yd��U���u�<�u�4��4�(���&���G��d��U���u�u�u�4��4�(�������@��Q��F��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��A���8�f�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʷ�:�
��,�"��O���&����CT�
N��Wʢ�0�u� �&�0�8�_����ԓ�l ��_�����i� �&�2�2�u��������EW��^�\���9�0�w�w�]�}�W���&����e9��h_�*��i�u�'�2��;�(��&���F��@ ��U��n�u�u�3���2���+����lU��^ �����3�
�a�
�e�a�W��Y����N��D�����8�
�b�3��n�(��Y�ƹ�@��R
�����;�!�9�d��m�F�������V�=N��U�������#�/�(�������T��B1�L���u�h�w�w� �8�Wǫ�
����WN��h��7���!�a�
�0��n�^������]��V�����
�#�f�d�g�t�W�������l�N��*���-� �
�l�1��@ׁ�H���U5��r)�� ���l�;�2�3��j�(��s���U5��r)�� ���l�;�2�3��j�(��E����`9��p����
�:�<�!�1��Aׁ�HӞ����T�����f�
�e�e�g�m�L���YӀ��}#��x��Dӊ�:�<�!�3��k�(��E�ƪ�l5��r-�� ���`�'�2�m�l�}�Wϸ�&����|��[�� ��l�%�u�h�1��2�������l��h��A���%�n�u�u�1��2�������l��h��A���%�u�h�}���0�������G	��Y�� ��l�%�u�:�w�-��������9��^�E���_�u�u����8���Jƹ��l��h��A���%�u�h�3���2�������l��h��D���%�n�u�u�1��2���-����S��h��A���%�u�h�_�w�}�W���*����K)��h_�����b�
�d�"�2�}����Kƹ��T9��F�U���d�|�0�&�w�}�W���YӀ��`#��t:����
�0�
�m�]�}�W���*����g)��h]��G���
�e�
�f�k�}�W���Y����`9��{+��:���f�
�=�
�"�l�B���Y����N��X��9��� �
�m�'�0�h�C��Y���O��[�����u�u�u����8���Jƹ��lR��h����u�x�u����4�������C��Q��Eߊ�a�4�&�2�w�/����W���F�Q=��0���� �
�d�'�4����Iƹ��l��^	�����u�u�'�6�$�u����O���� ��~ ��-���!�'�
�d�>�/��������R�Q=��0���� �
�d�%�:�F��Y����Z��D��&���!�
�&�
�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��P1������&�a�3�:�n�W���Y������T�����d�e�h�3���2���+����lR��^ �����'�2�`�a�~�t����Y���F�N��U�������#�n�(���&����S��N�U���'�c�$�n�w�}�W�������9F�N��U���u��������&����U��[��A��u��������&����V��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���-�
��-�"��D�������9��R�����9�2�6�#�4�2�_���������T�����d�
�|�x�"�.����Q����_T��h��*��|�n�u�u�>�8�(�������l��S��*���<�;�3�
�f��F�ԜY�ƥ�]��Q��Gߊ�f�i�u�'�0�����HĹ��P��S�����f�n�_�u�w�p����&Ź��W��D^�����;�%�:�0�$�}�Z���YӍ��A9��V
�����
�&�<�;�'�2�W�������@N��h��*���$��
�!��.�(������T9��R��!���f�3�8�g�w�0�(�������9��N����
� �a�a�'�t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���>�'�
�
�3�/���E�Ƹ�C9��h��A���%�}�f�x�f�9� ���Y����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�>�'�
��9����I���G��V�� ��a�%�}�f�z�l��������l�N��Uʰ�&�u�u�u�w�}�W�������9��S�����h�w�����/���[���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����
�
�0�u�$�4�Ϯ�����F�=N��U���'�c�6�e�6�.���������T��]���6�y�4�
�>�����*����9��Z1�U���&�2�6�0��	��������l�N�����u�u�u�u�>�}�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���K����lW���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�}����s���F�N�����
�
�0�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���X��hX�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F���*���
� �d�f�'�}�Jϭ�����Z��R�� �&�2�0�}�'�>��������O������1�%��&�;��(���H�ߓ�O�=N��U���0� �!�&�1��Bց�H���@��[�����6�:�}�0�>�8��������G��Q��@ۊ�f�y�a�|�]�}�W����ԓ�l ��X�����h�_�u�u�w�}����&¹��lW��h����u�<�;�2�1��Eځ�J���F�G�����_�u�u�u�w���������F9��1��N���u�%��9�����N����[�N��U���!�%�g�
�"�o�F���Y����N��G1�����g�
�g�e�w�}�F�������9F�N��U���
� �g�`�'�f�W���	����9��Q��Gۊ�g�i�u�!��2����������^	��¡�%�d�
� �d�j����Rӓ��Z��SF��#���
�
� �g�`�-�^��Y����l0��1�����l�
�f�i�w�}�W���YӒ��lT��Q��Bي�d�"�0�u�$�1����&����S��F�U���d�|�0�&�w�}�W���Yӕ��l��1��*��
�f�_�u�w�����O����W��G]��H�ߊu�u�u�u�/��2�������l0��B1�B���u�=�;�}�:��B�������V�
N��R���9�0�_�u�w�}�W����ԓ�l��h[�N���u�%�&�3��h�(��E��ƹF�N�����;�!�9�d���1ϩ�����@��h��D���%�}�|�h�p�z�W������F�N��*���&�
�#�a�g�W�W������� V��G]��H�ߊu�u�u�u�$�8�(���H�ӓ� F��R �����d�
� �g�b�-�_���D����F��D��U���u�u�!�%�e����H����9F���*���!�3�
�g��o�K�������T��A�����;�<�;�1�6�����&����lV�N�����0�}�8�
�a�;�(��&���l�N�����%�f�1�8�%�<�(���J�Փ�F�F�����%�
�0�:�0�3����MĹ��	��C��F���
�m�
�g�l�}�Wϭ�����9��h]�*��i�u�!�%�f�;�(��&����\��G1�����9�d�d�n�w�}��������U��]��G��u�!�%�c�1��Fց�KӇ����h��D���
�g�
�g�l�}�Wϭ����� 9��h]�*��i�u�u�u�w�}����K¹��lT��h����u�&�9�!�'����J����O�I�\ʰ�&�u�u�u�w�}��������_��h^�U���&�9�!�%��(�D���	���N��G1�����f�
�g�4�3�.����	���� Q��G\����u�0�
�8�a�9��������lU��h�I���!�%�d�3��j�(���Ƹ�C9��Q��Dӊ�g�n�u�u�$�1����&����U��N�U¦�9�!�%�
�2�2��������9����U���6�;�!�9�f�l�L���Yӕ��l�� 1��*���
�g�i�u�#�-�D���&����CT��Y
�����8�c�3�
�b��E��Y����V
��Z�����c�
�f�i�w�}�W���YӖ��R
��1��*��
�g�"�0�w�.����	Ĺ��lU��h�E���u�d�|�0�$�}�W���Y����V
��Z�����f�
�f�_�w�}��������lU��h�I���&�9�!�%�d�9��������lU��h����4�
�:�&��+�(���s���F�D�����4�!�3�
�f��F��Y����_	��T1�����}�0�<�0�$�:��������l ��^�����f�|�n�_�w�}��������V��G]��H�ߊu�u�u�u�:��(���H�ӓ�F��R �����f�3�
�m��o�G���Y�����RNךU���u�u�8�
��(�E���	��ƹF��Z��E���
�a�
�g�k�}��������E��X�����
�<�=�}�>�3�Ǯ�/����9��h_�*��y�:�<�!�0�/��������V�N�����3�
�a�
�f�n�Z�������V�G����u�u�u�8��l����O����Z�D�����6�#�6�:��8����
����WN��G1�*���g�`�%�|�d�t�L�ԜY�Ƹ�C9��h��G���%�u�h�&�3�1��������AN��^�����}�;�<�;�3�)���&����U��G�����!�2�'� �$�:����I���@��Z�����3�
�d�
�f�n�Z�������V�G����u�8�
�f�1��Oځ�K���W�@��U¦�2�0�}�8�����L����X��^	��´�
�:�&�
�!�o�D���Y����D��d��Uʡ�%�d�
� �f�j����Dӏ��T9��Q��D݊�d�`�u�u�w�2����I��ƹF��Z��@���
�l�
�g�k�}��������E��X�����1�4�
�:�$�����?���F��P ��]���3�
�m�
�e�t�}���Y����P��B1�B���u�h�&�1�;�:��������A��M�����;�1�$�
�"�n�N���P����]ǻN�����b�3�
�f��n�K���Y���F��Z��C���
�g�
�d� �8�WǼ�����v��C1�*���a�m�%�}�~�`�P���Y����l�N��Uʧ��6�&�
�"�i�O���B�����h_�����`�
�d�i�w�)�(�������P������� �&�2�0��0�(�������9��B�\��u�u�u�u�#�-�Fց�����F9�� 1��U��&�1�9�2�4�+����Q����I��^	��¡�%�d�
� �e�l����J���9l�N����
� �a�a�'�}�Jϭ�����Z��R��§�&�/�}�;�>�3�ǫ�&����J)��hZ�����`�l�y�a�~�W�W�������U�� Y��G��u�d�u�=�9�u����&����W��N�����:�&�
�#�d�m�W�������l�N����
� �g�`�'�}�JϮ�/����9��h_�*��d�u�u�u�8�3���B�����h\�����`�
�d�i�w�0�(�������9��_�X��1�"�!�u�~�W�W�������l ��Y�����h�!�%�d��(�E���	����K�
�����e�n�u�u�#�-�Eہ�����l��S��*���g�g�3�
�a��DǪ�&����T��B �����}�8�
�l�4�.�(���K�ѓ�O�S�����:�<�!�2�%�(�����θ�C9��h�����
�l�
�d�~�}����Q����]��R�����;�1�!�%�f���������9��G�U���;�u�:�<�#�:�ǫ�
����WN��G1�*���!�3�
�l��l�^��J�Ʃ�@�L�U���!�%�g�
�"�i�C���Y����l0��1�����d�
�f�d�w�}�W������]ǻN�����
� �g�d�'�}�Jϭ�����Z��R��§�&�/�}�;�>�3�ǭ�&����P��h��G���%�|�`�|�l�}�WϪ�	�Փ�F9��1��U��w�w�"�0�w�.����Q�ԓ�F9��1��\��&�2�0�}�'�>��������wO�R��U��n�u�u�!�'�i����@ƹ��Z�D�����6�#�6�:��4��������]��[�*���|�~�&�2�2�u�E���&����CT�d��Uʡ�%�`�3�
�g��E��Y����_	��T1�����}�;�<�;�3�<�(���
����T��N� ���2�0�}�g�1��O܁�K����F�C��C���
�d�
�g�k�}�F������uT��B1�F���u�u�%�6�9�)���&����_��^�����u�8�
�
�"�l�F���Y����A��a1��*��
�d�c�u�w�}�������9F���*Ҋ� �g�l�%�w�`�U���������^	��¦�
�8�
� �e�j����Eӓ��Z��SF��*���&�
�#�g�d�t�W�������l�N�����3�
�a�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���&����e9��h_�*��y�g�|�_�w�}��������l��S�����:�&�
�#��}�W���&�ғ�F9�� 1��\�ߊu�u�8�
��(�E���	���D�������;�<�;�1�$���������l��R�����;�1�4�
�8�.�(���K�����RN��W�ߊu�u��-��$����J����R��G\��Hʦ�1�9�2�6�!�>����������T�����d�
�e�e�w�}����ے��lW��Q��Fފ�f�|�_�;�w�8���