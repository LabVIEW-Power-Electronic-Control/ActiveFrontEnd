-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��A���Hŀ��l ��S����;�
�g�&�d��(���������N�����'�6�}�u�w�}�Wϗ�Y���F�N�����'�o�u�m�]�}�W���Y����`2��rN��U���0�0�u�h�d�W�W���Y�ƨ�]V��~*��U���;�0�0�u�j�n�L���Y�����1��1���o�<�!�2�%�g�W��s���F�S��*����u�u�;�2�8�W��J���F�=N��U���!�}�u�u�w�}����Y����Z�D�����6�_�u�u�w�}����Y����]F��C
�����n�u�u�u�w�>�W���Y�ƥ�F��S1�����_�u�u�u�w�4�G���Cӏ����h�����0�!�'�1�9��>���T�ƨ�D��^����u�u�u�<�f�}�MϷ�Yӕ��l
��^�����'�1�;�
��	�Z�������V�=N��U���u�%�:�0�m�4�Wϭ�����Z��R����1�"�!�u�~�W�W���Y�ƨ�F�T�� ���!�
�:�<��8��������d/��C����!�u�|�u�w�t�}���Y����G��=�����6� �0�4�4�}�ϳ�?����P��1����� �
�g�&�d�3�(���J����_9��GN�����u�x�x�x�z�p�Z��T���F��Z�����x�x�x�x�z�p�Z��T���9F������;�u��c�g�l��������W��B��*���9�1�%�f�w�.�W���Y����\��d��U���u�u�u�4�;�}�W���Y���F�N��U���;�u�!�
�8�4�L���Y���F������u�u�u�u�w�}�W���Y�ƥ�F��S1�����_�u�u�u�w�}�W�������l��[��U���u�u�o�<�w�.��������F�N��U���&�4�<�
��9����Y���F���U���
�:�<�
�2�)���Y����G	�UךU���u�u�u�u��%��������WF�N��U��<�u�&�1�;�:��ԜY���F�N�����
�
�1�!�w�}�W���Y����]F��C
�����
�0�!�'�d�}�������9F�N��U���u�
�-�&�8�8��������_��N��Uʦ�1�9�2�6�]�}�W���Y���@9��^�����!�:�
�1�#�}�MϷ�Yӕ��l
��^�����'�b�1�"�#�}�^�ԜY���F�N�����
�0� �!�#�<����Y����F��C
�����n�u�u�u�w�}�Wϳ�����A��[�����u�u�u�u�"�}��������E��X��Dʱ�"�!�u�|�w�}�W���P���F��SN�����0�!�_�u�w�p�Z��T���K�C�Xʙ�6�9�&�2�6�}�Z��T���K�C����u�<�;�9�6�1�W���Y�����h����u�u�&�2�6�}�������F��D�����6�_�u�u�>�3�Ͽ�����WF�T�����:�<�n�u�w�.����Y����R��N��Oʦ�1�9�2�6�!�>����Hӂ��]��G�U���&�2�4�u��+����Y����@��[���ߊu�u�<�;�;�?�������\��C
�����
�0�!�'�d�}�������9F������:�
�#�9�3�}�Mϭ�����Z��N�����4�u�%�!�6�<�W���Y����_	��T1�����}�u�:�;�8�m�L���Yӕ��]��E1�����u�u�o�&�3�1����s���@��V��*���!�u�u�u�w�)�(�������P��]����!�u�|�_�w�}����ӂ��9��Q_��U���!�
�:�<��8��������d/��C����!�u�|�_�w�}����ӂ��9��Q_��U���!�
�:�<��8��������d/��C����!�u�|�_�w�}����Ӊ��\��U��U���!�
�:�<��8����Hӂ��]��G����;�u�u�x�z�p�Z��T���K�C�����;�<�!�:�w�p�Z��T���K�d��Uʸ��a��c����������Q9��Q��*���
�g� �o�4�0����Ӌ��R��X��E���
�4�1�&�5�l����&���� TǻN�����8�%�}�u�w�}�WϿ����F�N��U���u�u�u�k�6�1�[���Y�����\��U���u�u�u�u�w�}�W�������]JǻN��U���
�-�&�4�#�<����Y���F������1�_�u�u�w�}�(���
����W��N��U���u�h�u�
�3�)�[���Y�����O�����4�<�u�u�w�}�W�������_��=N��U���u�
�-�&�5�)����Y���F�
P��*���!�y�u�u�w�}��������V��^�����<�u�k�:��+����s���F�D1�����%�'�!�:��9����D�ƣ�l��C�U���u�u�8�4�>���������_��N��Kʧ�!�4�<�y�w�}�W�������@9��D��*���!�u�u�u�i�/�������O��=N��U���x�x�x�x�z�p�Z��T�ƍ�@��Z��U���x�x�x�x�z�p�Z��T�����\N��U���h�6�>�_�w�}�������[��RUךU���
�#�9�1�w�`�P���s���R9��V��U��u�1�;�
��	�Z�������V�	N��R���=�;�}�1�9����D����Z��`'��=��1�"�!�u�w�c�P���P�ƣ�N��Y^�� ��h�}�1�;���#��Y����G	�S�R��|�u�9�0�3�3�(���H���F��C�����i�u�d�n�w�}�������Z�
��D�����d�1� �)�W���G����F��R ��]���d�7�3�u�w�}����.����W��X����h�u��|�w�2�WǺ�¹��UW�F��������d�3�*����Y���fA�N�����<�d�7�3�l�}�Wϱ�&����Z�
N��R�ߊu�u�%�!�6�<�W��[����V��N�����}�%�:�0�5�;�W���!���\�X����� �d�h�w��t�W������V��^��Sʺ�6�1�
� �f�f�W�������F�R�����4�4�_�u�w�p�Z��T���K�C�X���;� �u� �1�/�Z��T���K�C�X���u�%�:�0�$�u��������9F�N��U���6�>�0�0�#�<�Ͻ����A��_��U���u�u�u�u�>�}���^����[��N��U���u�u�u�u�3�3�(���H���F��Y^�U���u�u�u�u�w�}����&����F�
N����u�u�u�u�w�}�W�������V9��Q_��Hʺ�6�1�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��ʴ�6�<�0�!�%�f�