-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�g�e�f����(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�4�0��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�^ �����
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W�������T��h��U���������!���6���F��@ ��U���_�u�u�;��3�������/��d:��9�������w�n�W������]ǻN�����;�0�b�0�c�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��a��R1�����o��u����>���<����N��
�����e�n�u�u�>�����&Ĺ��F��~ ��!�����
����_������\F��d��Uʼ�
�4�2�
���W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V �����!�:�
�g�2�m�Mϗ�Y����)��tUךU���;��;�4��3����H����F��~ ��!�����
����_������\F��d��Uʼ�
�4� �9�8�)����K����\��yN��1�����_�u�w�3�:�������G��h_����o��u����>���<����N��
�����e�n�u�u�>���������A	��\��*���u������4�ԜY�ƥ�l+��B�����:�
�g�0�b�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��~��V�����9�d�
�
�w�}�9ύ�=����z%��N�����4� �9�:�#�2�(������/��d:��9�������w�n�W������]ǻN�����<�&�a�0�g�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Yӏ��t��D1����o��u����>���<����N��
�����e�n�u�u�>�����&ǹ��F��~ ��!�����
����_������\F��d��Uʼ�
�4�;�
���W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V��*ފ�
�u�u����;���:����g)��]����!�u�|�_�w�}��������l��T��;ʆ�������8���J�ƨ�D��^����u�;��<�$�i���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF��Y1�����a�0�b�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϷ�&����G9��N��U���
���n�w�}����/�ԓ�lV�'��&���������W��Y����G	�UךU���;��
�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƥ�l6��1��G���u��
���(���-��� W��X����n�u�u�<���E���J����}F��s1��2������u�d�}�������9F���&���
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���*����V9��N��U���
���
��	�%���Hӂ��]��G�U���4�
�0� �9�m�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���R��R����o������0���/����aF�N�����u�|�_�u�w�-��������	F��cN��1��������}�D�������V�=N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӇ��A��E ��U��� �u��
���(���-��� W��X����n�u�u�4��8����L����f2��c*��:���
�����l��������l�N��*��� �;�c�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���	����F�� N�:���������4���Y����W	��C��\�ߊu�u�%�'�#�/�(���Y����`2��{!��6�����u�f�w�2����I��ƹF��G1�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}��������}F��s1��2���|�_�;�n�]�<��������VF��_�����e��c�a�1�m�����ƹF��X �����4�
�:�&��2����Y�Ɵ�w9��p'��O���d�n�u�u�4�3����Y����\��h�����u�u��
���W��^����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�g�u�8�3���Y���V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�
�&��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�d�w�]�}�W���
������d:��ي�&�
�u�u���8���&����|4�]�����:�e�u�h�u�m�G��I����V��^�E��w�_�u�u�8�.��������l��h��*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
�ӓ�@��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��H����]ǻN�����4�!�4�
��.�A������5��h"��<������}�d�9� ���Y���F�^�E��e�e�e�e�g�m�G��B�����D��ʴ�
��&�b�1�0�A��*����|!��h8��!���}�f�1�"�#�}�^��Y����V��^�E��e�d�e�e�g�f�W�������R��V��!���m�3�8�b�m��3���>����v%��eN��Fʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�����m�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W���*����V��D��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6��#���H¹��^9��T��!�����
����_������\F��T��W��e�e�e�e�g�l�G��I����]ǻN�����4�!�4�
��.�F݁�
����\��c*��:���
�����n��������\�^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
��&�f�����K����g"��x)��*�����}�f�3�*����P���V��^�E��d�e�e�e�g�m�G��Y����\��V ������&�d�
�$��D��*����|!��h8��!���}�f�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�f�W�������R��V��!���d�
�&�
�c�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�n�w�}��������R��c1��D܊�&�
�`�o���;���:����g)��\����!�u�|�o�w�m�G��I����V��^�E��e�n�u�u�4�3����Y����g9��Y�����c�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W���*����^��D��B��������4���Y����W	��C��\��u�e�e�e�f�m�G��I����V��L�U���6�;�!�;�w�-�$����ߓ�@��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����D��N�����!�;�u�%����������
F��d:��9�������w�o�W������F��L�E��e�e�e�e�g�m�G��I����F�T�����u�%��
�#�l����K����`2��{!��6�����u�g�w�2����I����D��_�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�g�1�0�E���Y����)��t1��6���u�g�u�:�9�2�G���D����V��^�E��e�e�e�e�g��}���Y����G����&���!�f�3�8�e�}�W���&����p9��t:��U��u�:�;�:�g�}�J���H����V��^�E��e�e�e�w�]�}�W���
������d:�����3�8�g�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y�����d�o�����4���:����V��X����u�h�w�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�d�e�u�W�W�������]��G1�����9�f�
�e�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�d�g�m�L���YӅ��@��CN��*���&�
�#�g��g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�l�F��Y����\��V �����:�&�
�#�e�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���e�1�"�!�w�t�M���I��ƹF��X �����4�
�:�&��+�E��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$�����J����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����W��UךU���:�&�4�!�6�����&����lP�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h_�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��A]��D���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��d�w�_�u�w�2����Ӈ��P	��C1��F؊�a�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�d�e�n�w�}��������R��X ��*���g�d�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�f�
�c�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�d�f�m�L���YӅ��@��CN��*���&�
�#�g�f�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d�m�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����F�T�����u�%�6�;�#�1�E��Cӵ��l*��~-��0����}�u�:�9�2�G���D����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�d�3�*����P���W��d��Uʶ�;�!�;�u�'�>�����ԓ�\��c*��:���
�����}�������	[�^�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��_�W�ߊu�u�:�&�6�)��������_��h/��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[��A��������4���Y����\��XN�U��w�e�w�_�w�}��������C9��Y�����d�o�����4���:����T��X����u�h�w�e�u�W�W�������]��G1�����9�f�
��m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�d�f�m�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Bʱ�"�!�u�|�m�}�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�g�w�2����I����D��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#�b�i�G���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�n�u�u�4�3����Y����\��h��@��e�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����D��N�����!�;�u�%�4�3����A����	F��s1��2������u�`�9� ���Y���F�_�D��n�u�u�6�9�)����	����@��A_��@��o������!���6���F��@ ��U���o�u�e�e�f�l�G��I���9F������!�4�
�:�$�����H���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����d�
�e�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��L�U���6�;�!�;�w�-��������9��N��1��������}�NϺ�����O�
N��E��e�e�e�n�w�}��������R��X ��*���m�f���m��3���>����v%��eN��Bʱ�"�!�u�|�m�}�F��H����W��_�D��u�u�6�;�#�3�W�������l
��1��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�F��H���9F������!�4�
�:�$�����H����g"��x)��*�����}�b�3�*����P���V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�g�b��g�m�W���-����t/��a+��:���f�u�:�;�8�m�W��[����W��_�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����F��d:��9�������w�i��������\�^�E���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Mӂ��]��G��H���e�e�w�_�w�}��������C9��Y�����a�o�����4���:����R��X����u�h�w�e�g��}���Y����G�������!�9�`�g�m��3���>����v%��eN��U���;�:�e�u�j��G��[��ƹF��^	��ʴ�
��3�8�m��3���>����v%��eN��Fʱ�"�!�u�|�m�}�G��I����V��^�E��e�d�n�u�w�<��������@��Y�����o�&�'�;�l�}�WϿ�����G��D�����<�2�:�u�'��(���Y�ƿ�T����W���0�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��o�MϜ�6����l�N�����u�'�
����<���	����Q��B����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����u#��u/����� �
�d�
�"�;���Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������4�'������������9��Q��*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4��������v#��v-�� ���!�g�b�7�1�8�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����'�
������������l��Q��C��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:��������v"��t%�����
�d�
� �1�/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʴ�'�����2����&����Q��R��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�>�3�Ͽ�����w$��|�����g�b�7�3�2��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��P ��U���
�����(����Aƹ��	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�'���3���2����F��1�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�&�0�<�W���&����
W��N�&���������W��Y����G	�UךU���<�;�9�'�0�l�F���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�D�������	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��R��!���d�
�&�
�a�g�$���5����l�N�����u�%�&�2�5�9�F��CӤ��#��d��Uʦ�2�4�u�'��(�N���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʧ�2�d�g�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�l��h�����
�!�a�3�:�l�W���-����t/��=N��U���;�9�4�
�>�����K����q)��r/�����u�<�;�9�>�����&ù��R��R�����d�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����u#��u/����� �
�d�
�"�;��������
R��N��1��������}�D�������V�=N��U���;�9�4�'���5�������G9�� 1�����
�
�0�
�n�e�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��0����� �%�#�o�@�������9��P1�@���u��
����2���+������Y��E��u�u�&�2�6�}����<����p-��C��*��
� �3�'�d�/���L����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�'�����2����&����Q��R��*���
�l�f�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��l ��s,��>���%�!�g�b�5�;����&����_��T��!�����
����_������\F��d��Uʦ�2�4�u�'���3���2����F��Y�� ���'�c�'�2�e�j�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V��3�����:�!�"��F؁�����lQ��R	��L��o������!���6���F��@ ��U���_�u�u�<�9�1��������P��N�&���������W������\F��d��Uʦ�2�4�u�
��8�(��O����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$���݁�
����	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������9��h_�G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����@ǹ��T9��_��U���
���
��	�%���Y����G	�UךU���<�;�9�0�>�>��������V��N�&���������W������\F��d��Uʦ�2�4�u�'���3���2����F��1�����
�0�
�l�o�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h(��1���� �%�!�o��(�������lU��N�&���������W��Y����G	�UךU���<�;�9�&�;�)����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�����I���5��h"��<������}�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��Z�Oʗ����_�w�}����ӕ��l��1��*��b�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��E��F��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������U��_�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	ǹ��T9��_��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%��2���:����C��_��F���e�g�3�
�f�h����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��������:�#�(�(��&����9��E��F��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����q'��X�� ���d�
�
�
�����Jʹ��\��c*��:���
�����l��������l�N�����u�'�
����<���	����Q��h��*ߊ�0�
�e�a�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��r+��4��� �%�!�g�`�n����A����W��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�/�1���;����F��C1�B���0�e�m�'�0�n�D���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��������:�#�(�(��&����9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������v#��v-�� ���!�g�b�f�2�m�Fށ�����R�=��*����
����u�FϺ�����O��N�����4�u�'�
���6�������lT��h]��*ۊ�
� �d�m��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��G1�����0�
��&�c�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}����<����p-��C��*��
�
�
�
��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����'�
������������lU��h_��*���d�g�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��r+��4��� �%�!�g�`�n����H¹��lW�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(�������^9��1��D���
�g�e�%�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�`�3�:�i�Mύ�=����z%��N�����4�u�%�&�0�?���H����|)��v �U���&�2�4�u�%���������W��1�����g�g�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ʃ�Z��Y
�����g�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l��R1�����d�
�
�
�"�l�@߁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
� �d�m��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��*���$��
�!��.�(���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<����<����x	��G��G���0�e�f�f�1��D���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʰ�<�6�;�f�1��E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�����(����K�ѓ�lV��h]�� ��`�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��l ��s,��>���%�!�g�b�2�m�F�������^��N�&���������W��Y����G	�UךU���<�;�9�4�%��2���:����C��_�����e�f�3�
�d�k����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��������:�#�(�(��&���� 9��Q��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������v"��t%�����
�d�
�
���(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�'�
���6�������lT��h��*ۊ�
� �d�a��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��0����� �%�#�o�@���H�֓�l ��Z�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l*��G1�*���d�c�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƥ�l
��q��9���
�c�'�2�d�n�W���-����t/��a+��:���g�1�"�!�w�t�}���Y����R
��G1�����0�
��&�`�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������U��Y�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�Г�V��Z�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�/�)����&����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������P��N�&���������W������\F��d��Uʦ�2�4�u�0��0�F؁�����T�=��*����
����u�W������]ǻN�����9�&�9�!�'�e����L�֓�F��d:��9�������w�m��������l�N�����u�0�
�8�f�����H���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�����2����&���� 9��1�*���d�e�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��r+��4��� �%�!�g�`�n����Hƹ��T9��^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��2���8����G��h\�*ي�
�
�`�3��h�G���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y���������8�)����HĹ��V9��[�����g�e�o����0���/����aF�N�����u�|�_�u�w�4��������l ��h"����
�
�
� �f�h�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�:�
�:�'�o�(���&���� T��T��!�����
����_������\F��d��Uʦ�2�4�u�9�;���������9��1��*���d�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��E1�����`�0�d�'�0�n�E���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����'��:��j��������
W��N�&���������W��Y����G	�UךU���<�;�9�6��)�1���5����Q��h^�����g�b�o����0���/����aF�N�����u�|�_�u�w�4��������l ��h"����
�
�
� �f�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�:�
�:�'�o�(���&���� T��T��!�����
����_������\F��d��Uʦ�2�4�u��;���������9��h_�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������A9��X��D���2�f�a�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l
��q��9���
�f�3�
�a�n����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����'��:��n����J����	F��s1��2������u�d�}�������9F������6�
�!��%�����L����l ��X�*��o������!���6�����Y��E��u�u�&�2�6�}����&����	��h]�����'�2�f�`�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������_9��h(��*���%�f�
�
��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����9�9�
�:��2���&����A��\�U����
�����#���Q����\��XN�N���u�&�2�4�w����� ����S��R	��G��o������!���6���F��@ ��U���_�u�u�<�9�1��������V��c1��Dڊ�&�
�u�u���8���B�����Y�����<�
�1�
�a�}�W���5����9F������3�
���e����&����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����-����G9��h\�����g�c�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����O����T9��_��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�1�(���&����lT��1��E���3�
�l�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�g���(߁�&���� T��T��!�����
����_������\F��d��Uʦ�2�4�u�%�$�:����&����GW��Q��D���u��
���f�W���
����_F��h��*���
�m�u�u���6��Y����Z��[N�����
�:�
�:�'�o�(܁�&ù��U��_�����u��
����2���+������Y��E��u�u�&�2�6�}��������l*��G1�*ي�
�
�
�0��o�F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*����'��:��e�D���I�ѓ�F9��[��F��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h\��F���e�b�'�2�d�d�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e��(���&�֓�F9��X��F��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h\��F���e�d�
�0��n�F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*����'��:��e�D���H�ד�F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h\��F���d�d�'�2�d�m�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e��(���&ǹ��lW�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���?����\	��V��*���
�
�0�
�d�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�o�n����N����_��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�/��������\��1�����b�'�2�f�f�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�g���(ށ�I����V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�/��������\��1�����d�
�0�
�d�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1��9����!�`�
�"�o�Eف�J����g"��x)��*�����}�d�3�*����P���F��P ��U�������#�h�(���&����\��c*��:���
�����l��������l�N�����u�%�&�2�4�8�(���
����U��W��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��G1�*���g�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��*��b�o�����4���:����V��X����n�u�u�&�0�<�W���
����@��d:�����3�8�g�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��l�W���6����}]ǻN�����9�!�%�m��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�m�
�0��n�E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����d�<�3�
�e�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
�
�0��n�O��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����e�<�3�
�e�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
�
�0��n�C��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����l�<�3�
�e�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
�
�0��n�G��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����b�<�3�
�e�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���f�
�
�0��n�A��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e��(ށ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�%�$�:����&����GT��Q��G���u��
���f�W���
����_F��h��*���
�f�u�u���6��Y����Z��[N�����
�:�
�:�'�o�(܁�&���� _��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%���������C9��h]��*���g�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��C1�����:�
�g�f�f����Jǹ��\��c*��:���
�����l��������l�N�����u�'�
�!��/�;���&�Г�l��h_�� ��a�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��l
��q��9���
�c�f�0�g�i����M�ӓ� F��d:��9�������w�n�W������]ǻN�����9�4�'�9��2�(���	���� 9��1�����a�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�A9��h(��*���%�f�
�
���F���&����l��N��1��������}�D�������V�=N��U���;�9�4�'�;���������9��R1��D���
�`�a�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��[�����:�%�f�
���(ہ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��)�1���5���� P��h��*݊� �g�f�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��3����:�
�c�d�8�F��&����S��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�����Oʹ��\��c*��:���
�����}�������9F������4�
�<�
�$�,�$����Փ�@��N�&������_�w�}����Ӈ��@��U
��A��o�����W�W���������h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:����	����l��F1��*���a�3�8�g�w�}�#���6����9F������4�
�<�
�3��@���Y����v'��=N��U���;�9�4�'���5�������G9�� 1��D���'�2�f�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��r+��4��� �%�!�g�`�8�F�������R�=��*����
����u�FϺ�����O��N�����4�u�'�
���6�������lT��h]��*ۊ�
�0�
�m�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��q+��7���:�!� �
�f��(���&ʹ��T9��N�&���������W��Y����G	�UךU���<�;�9�4�%��2���:����C��_�����f�'�2�a�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h(��1���� �%�!�e�j����K����lR��T��!�����
����_������\F��d��Uʦ�2�4�u�'���3���2����F��Y��*���
�
�0�
�d�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��E1��0����:�!� ��l�(܁�&ù��A��Z�Oʆ�������8���J�ƨ�D��^����u�<�;�9�>�/���A����g"��x)��*�����}�u�8�3���B�����Y���������8�)����HĹ��V9��E��A��o������!���6���F��@ ��U���_�u�u�<�9�1����?����r%��B����b�e�0�d�%�:�C��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����:�0�!�'��l�(܁�&����_��N��1��������}�D�������V�=N��U���;�9�4�'�9�9�(�������lT��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����l��Z1�@���'�2�`�l�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�A9��r*��6���!� �
�d���(܁�&����U��N��1��������}�D�������V�=N��U���;�9�4�'���5�������G9�� 1��D���g�'�2�`�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h(��1���� �%�!�e�j����H�ԓ�V��^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��2���8����G��h\�*���
�
�
�0��k�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V��3�����:�!�"��F؁�&ù��9��P1�E��������4���Y����W	��C��\�ߊu�u�<�;�;�<����<����x	��G��G���0�e�g�g�%�:�B��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V���������"�-���N����lW��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����q'��X�� ���d�
�
�
������I����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʼ�
�0�
�d�w�}�#���6����e#��x<��Gʱ�"�!�u�|�]�}�W�������_9��s+��'���'�
�g�
������K����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʶ�
�����8���M����l��hX�U����
�����#���Q����\��XN�N���u�&�2�4�w�1�>���!����V��\�����'�2�c�`�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������_9��s+��'���'�
�g�
������L����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʶ�
�����8���O����l��hX�U����
�����#���Q����\��XN�N���u�&�2�4�w�1�>���!����V��\�����'�2�c�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������_9��s+��'���'�
�g�
������@����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʶ�
�����8���I����l��hY�U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(�������^9��h_�����d�u�u����>���<����N��
�����e�n�u�u�$�:��������W��R��Mۊ�
�0�
�g�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����P
��b ��0���8�d�l�0�g�/���H����g"��x)��*�����}�d�3�*����P���F��P ��U������!�%��@ց�&¹��T9��N�&���������W��Y����G	�UךU���<�;�9�6���3�������_��h^�����c�u�u����>���<����N��
�����e�n�u�u�$�:��������w*��R��D���0�g�'�2�`�j�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��[1��;���!�'�
�c���(���&����	F��s1��2������u�d�}�������9F������6�
� ���8���@����l��hV�U����
�����#���Q����\��XN�N���u�&�2�4�w�1�5���5����^9��1��D���2�m�f�o���;���:����g)��]����!�u�|�_�w�}����Ӆ��q3��{+�����c�
�
�
�2��E���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*�����0�8�f�d�������� Q�=��*����
����u�FϺ�����O��N�����4�u�9�������&����V9��E��M��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��X��C���0�e�'�2�o�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�a�n����K����l^��T��!�����
����_������\F��d��Uʦ�2�4�u�'��)�1���5���� P��h^��*���0�
�m�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�A9��h(��*���%�f�
�
���(���&����	F��s1��2������u�d�}�������9F������4�'�9�
�8�����JŹ��V9��E��L��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��X��C���0�d�g�'�0�d�F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*����'��:��k����K����V��]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%���������C9��h��*ي�
�0�
�a�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Z*��^1�����:�
�
�0��h�W���-����t/��a+��:���g�1�"�!�w�t�}���Y����R
��1����m�o�����4���:����T��X����n�u�u�&�0�<�W�������9��h\�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�܁�����
F��d:��9�������w�l��������l�N�����u�-�!�:�3�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����'�
�!��%�����O�Փ�lV��1��*��f�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����V��Q��@���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�����u	��{��*���f�0�d�d��(�E��&���5��h"��<������}�f�9� ���Y����F�D�����'�
�:�0�#�/�(�������C��Q��B���%�u�u����>���<����N��
�����e�n�u�u�$�:��������9��h\�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��(�N���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��V�Oʗ����_�w�}����Ӈ��@��T��*���&�d�
�&��m�Mύ�=����z%��N�����4�u�%�&�0�?���L����|)��v �U���&�2�4�u�'�.��������l��1����u�u��
���L���Yӕ��]��V�����1�
�e�u�w��;���B�����Y�����3�
�l�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��L���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l_��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-����@ʹ��\��c*��:���
�����l��������l�N�����u�8�
�g�1��G���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʡ�%�b�
� �f�m�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����`�3�
�e�`�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��Bߊ� �d�e�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hY�����e�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������v#��v-�� ���!�g�b�f�2�m����I�ߓ� F��d:��9�������w�n�W������]ǻN�����9�4�'����4�������W��1��E���3�
�d�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��E1��0����:�!� ��l�(܁�&ù��U��\�����u��
����2���+������Y��E��u�u�&�2�6�}����<����p-��C��*��
�
�
�
��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����'�
������������lU��h^��*���d�a�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��r+��4��� �%�!�g�`�n��������W��N�&���������W��Y����G	�UךU���<�;�9�4�%��2���:����C��_��F���d�d�3�
�f�e����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��������:�#�(�(��&����9��Q��D���%�u�u����>���<����N��
�����e�n�u�u�$�:��������v"��t%�����
�d�
�
���(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�'�
���6�������lT��h]��*ۊ�
� �d�d��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��@���
�g�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������\��Q��G���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�����V9��E��D؊�
� �d�`��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��C���
�g�e�%�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������V
��Z�����g�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1��*��m�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��Q��F���%�u�u����>���<����N��
�����e�n�u�u�$�:��������CW��B1�G؊�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l ��]�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������U��]�����u��
����2���+������Y��E��u�u�&�2�6�}�����ӓ�F9��Z��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�֓�F9��^��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�ד�F9��Z��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�ԓ�F9��\��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�Փ�F9��V��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�ғ�F9��X��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�ӓ�F9��\��F��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����P��G_��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%��2���:����C��_��F���e�d�
� �f�j�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V���������"�-���N�Փ�lV��1��*��g�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����u#��u/����� �
�d�
���(�������R��N�&���������W��Y����G	�UךU���<�;�9�4�%��2���:����C��_��F���d�d�
� �f�o�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�d�
� �f�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�i�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�h�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�j�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�e�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�d�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�m�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�o�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�g�
� �f�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�f�
� �f�i�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����8�f�
� �f�k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�d�3�
�a�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���f�
� �d�a��F��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����d�3�
�c�g�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��[1��*���
�:�%�f���(���H����CW�=��*����
����u�W������]ǻN�����9�&�9�!�'�o����O�Г� F��d:��9�������w�m��������l�N�����u�0�
�8�d����Aù��\��c*��:���
�����l��������l�N�����u�0�
�8�d����AŹ��\��c*��:���
�����l��������l�N�����u�� �������&�ԓ�F9��^��D��������4���Y����W	��C��\�ߊu�u�<�;�;�1��������U��N�&���������W������\F��d��Uʦ�2�4�u�:���E���&����l��N��1��������}�E�������V�=N��U���;�9�!�%�>�4���&����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�4��������Q��N�&���������W������\F��d��Uʦ�2�4�u�0���(�������
9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��n�(���&����lW�� 1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�%�)�E�������R��T��*���d�a�
�f�m��3���>����v%��eN��Aʱ�"�!�u�|�]�}�W�������V
��Z��*���d�`�
�f�m��3���>����v%��eN��Aʱ�"�!�u�|�]�}�W�������l4��B�����
�b�l�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����U5��z;��G���!�m�
�;�2�-�!�������Q��N�&���������W��Y����G	�UךU���<�;�9�!�'�4����N�Փ�F��d:��9�������w�m��������l�N�����u�8�
�d�����@ʹ��\��c*��:���
�����}�������9F������!�%�`�
�"�l�Gځ�K����g"��x)��*�����}�u�8�3���B�����Y�����c�
� �d�f��D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Lӊ� �d�g�
�f�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��_�� ��f�
�f�o���;���:����g)��Y�����:�e�n�u�w�.����Y����W��h�� ��d�
�f�o���;���:����g)��\����!�u�|�_�w�}����Ӓ��l^��^1��*��l�%�u�u���8���&����|4�^�����:�e�n�u�w�.����Y����@��hY�����m�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l��{:��:���m�
�;�3��-�(���H����CU�=��*����
����u�CϺ�����O��N�����4�u�0�
�:�k����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�j����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�e����&����l��N��1��������}�GϺ�����O��N�����4�u��-��	����&�ғ�F9��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;�3����&����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�1�(���&����lT��1��E���3�
�l�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�g���(߁�&����
T��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%���������C9��h]��*ڊ�
� �d�g��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�o�n����A����_��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�/��������\��1�����l�3�
�l�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e��(���&����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���?����\	��V��*���
�
� �d�o��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*����'��:��e�D���H�Г�F9��_��F��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h\��F���d�m�3�
�g�h����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�:�
�:�'�o�(܁�&¹��U��_�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K����U��]�����u��
����2���+������Y��E��u�u�&�2�6�}����&�Փ�F9��[��A��������4���Y����\��XN�N���u�&�2�4�w�2�(���M����V��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�O����V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�;�>�!��&����Q��GZ��U���
���
��	�%���Y����G	�UךU���<�;�9�9�4��Fف�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8���D���J����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�N����W��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�;�>�!��&����V��GZ��U���
���
��	�%���Y����G	�UךU���<�;�9�9�4��Fׁ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8���C���J����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�9�)��������U��N�&���������W������\F��d��Uʦ�2�4�u�:�;�.�(���K����CT�=��*����
����u�W������]ǻN�����9�;�!�=�a�;�(��H����	F��s1��2������u�g�9� ���Y����F�D�����:�9�&�
�"�o�Bځ�K����g"��x)��*�����}�u�8�3���B�����Y�����c�
� �g�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��C܊� �g�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��Y�� ��b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����U��W��G��������4���Y����\��XN�N���u�&�2�4�w�2����&����_��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�;�#�5�@���&����l��N��1��������}�GϺ�����O��N�����4�u�8�
�g�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����8�
�d�3��o�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����g�3�
�e�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@���
�e�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������W��R�����<�3�
�e�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��Gي�0�:�2�;�>�;�(��H����	F��s1��2������u�g�9� ���Y����F�D�����8�
� �g�d��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��D���1�8�'�4�����O¹��\��c*��:���
�����}�������9F������!�%�c�
�"�o�@ց�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�m�<�3�0����&����R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�j�(���K����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�e����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�(�������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�F�������F9��W��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������W��N�&���������W������\F��d��Uʦ�2�4�u�0��0�Eׁ�&����Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�k�(���K����CT�=��*����
����u�W������]ǻN�����9�!�%�b��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʳ�
����"��Gف�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�=�#�-����&����l��N��1��������}�D�������V�=N��U���;�9�&�9�#�-�E�������^��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������U��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�$�1����I����F9��^��F��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���¹��9��Q��F���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����^W��\��*���g�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V
��Z�*��� �g�`�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��@ڊ�
� �g�`��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��R�����
�
� �g�a��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����7����!�'�
�o�8�E���&����l��N��1��������}�D�������V�=N��U���;�9�4�'�;���������9��1��*��`�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����_��X�����g�
�
�
�"�o�Nց�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�!��'��2�(���J�Г�F9��X��F��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h\��F���3�
�a�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�g���(���K����CU�=��*����
����u�FϺ�����O��N�����4�u�����8���H�Г�l ��]�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��X��C���0�e�f�3��i�O���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�:�
�8�-�Dف�&����9��h\�G���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����\��X��F܊�
�
�
�
�"�o�Aց�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�!��'��2�(���J����l^��B1�Mي�f�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�����u	��{��*���f�0�e�l�1��C���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�'�9�
�:��2���&����9��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��h"����
�
�
�
��(�E��&���5��h"��<������}�f�9� ���Y����F�D�����'�
�!��%�����O�Փ�lW��h��G��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������G9��E1�����c�f�0�d�o�;�(��J����	F��s1��2������u�d�}�������9F������4�'�9�
�8�����JŹ��V9��1��*���l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G��1��*���l�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l ��h"����
�
�
�
�e�;�(��L����	F��s1��2������u�d�}�������9F������&�9�!�%�`�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����'�
�!��%�����O�Փ�lV��1��*���l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����_��X�����f�
�
�
��o����O�ӓ� F��d:��9�������w�n�W������]ǻN�����9�4�'�9��2�(���	���� 9��1�*���g�`�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��B1�D���6�1�u�u���8���&����|4�N�����u�|�_�u�w�4��������F9��1��U����
���l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����N���$��{+��N���u�&�2�4�w�-��������`2��C_�����d�u�u����>��Y����Z��[N��*���
�1�
�b�`�g�5���<����F�D�����%�&�2�6�2��#���HŹ��^9��T��!�����n�u�w�.����Y����Z��S
��B��o�����W�W���������D�����
��&�d��.�(��Cӵ��l*��~-�U���&�2�4�u�'�.��������F��u!��0���_�u�u�<�9�1��������
9��T��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�@݁����� 9��T��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�@ځ�����9��T��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�@ց�����9��T��U����
�����#���Q�ƨ�D��^����u�<�;�9�6��$�������g"��x)��*�����}�f�3�*����P���F��P ��U���&�2�7�1�e�i�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����R��N��:����_�u�u�>�3�Ͽ�&����Q��_�U������n�w�}�����ƭ�l��h��*��m�o�����}���Y����R
��G1�����1�g�a�u�w��;���B�����Y�����<�
�1�
�f�l�MϜ�6����l�N�����u�%�&�2�5�9�A��CӤ��#��d��Uʦ�2�4�u�%�$�:����K����	F��x"��;�ߊu�u�<�;�;�<�(���&����Q��N��:����_�u�u�>�3�Ͽ�&����Q��_�U������n�w�}�����ƭ�l��h��*��d�o�����}���Y����R
��G1�����1�g�c�u�w��;���B�����Y�����<�
�1�
�f�h�MϜ�6����l�N�����u�%�&�2�5�9�E��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߠu�u�6�8�8�8�ϳ�K���� ��1����� �
�g�&�d�3�(���J����_9��GN�����u�0�0�<�w�W�W���Y�ƅ�\��y:��0��u�u�u�u���$���<����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�<�d����Mϗ�-����l�N��Uʱ� �
���w�}�9���<���9F������u�u�u�u�4�6�Mϗ�Y����)��tUךU���u�u�0�0�w�}�9ύ�=����z%��N��U���1�;�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����\��yN��1��������}�D�������V�=N��U���u�%�:�0�m��W���&����p9��t:��U��1�"�!�u�~�W�W���Y�Ư�\��yN��1�����_�u�w�}�W�������f2��c*��:���
�����l��������O��N�����6�8�:�0�#�W�}���Y����\��CN��G��f��
�
�:�1�Dݰ�&�Ԣ�lU��1�����%��_�u�w�8����Y���F�N��U������n�w�}�W���7����g'��T��;����n�u�u�w�}����&����{F��~ ��2���_�u�u�u�w�4�F���=���/��r)��N���u�u�u�1�"��>���Y�ƅ�g#��eN����u�:�!�}�w�}�W�������	F��=��*����
����u�FϺ�����O��N��U���1�;�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����\��b:��!�����
����_������\F��G�U���0�1�6�8�8�8��Զs���P	��X ��ʸ�g�e�f�������J���� T��h_��U���u�u�2�;�%�>�_���Y���/��N��!����_�u�u�w�}�"���-����	F��c+��'�ߊu�u�u�u�>�m� ���1����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�:�!����Mϗ�-����O��N�����u�_�u�u�w�}���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N����o��u����>���<����N��
�����e�n�u�u�w�}��������z(��c*��:���
�����}�������9F�N��U���!�o�����;���:����g)��^�����:�e�u�n�w�}��������]��dװ���<�_�u�u������
������\��*���f�3�9�
�$��F���Y����\��CN��G��f��
�
�6�9����J���� T��h]��F���9�
�&�_�w�}�����ơ�CF�N��U����u�k�d�]�}�W���Y����`2��rN��U���u�u�u�u�3�3�(���-���U��=N��U���u�<�d����J���K���F�N�� �����u�k�d�t�W���	����^��d��U���u�6�>�h�w�-����s���F�E����u�%�'�!�]�}�W���Y����[�P�����l�
�e�_�w�}�W������F��G1��*��
�d�_�u�w�}�W������F��G1��*��
�%�:�0�]�}�W���Y���F��G1��*��
�0�_�u�w�}�W������T��Q��Lۊ�g�n�_�u�w��(�������@9��Y��G���8�-�1�%��m�MϽ�����]��\��C���3�e�3� ��o�������lW��V���ߊu�u�0�0�>�}����s���F�~*��K��_�u�u�u�w��(���>���W�N��U���1�;�
���}�I��U���F�
��D�����h�u�e�W�W���Y�ƨ�F��~*��U��f�|�u�u�'�/�W���Y���F�N�����k�2�%�3��d�(��s���F�S��U��2�%�3�
�n��F�ԜY���F��B��Kʲ�%�3�
�l��o�L�ԜY�ƪ�9��Z��G���f�;�
�
��o�W�������V��Z^��E���
�
�6�'�n����K����lWǻN�����<�u�4�u�]�}�W���Y���F��=N��U���u� �
���}�I��s���F�S��*����u�k�f�{�}�W���Yӂ��9��s:��H���g�_�u�u�w�}����.����[�GךU���:�!�8�%��}�W���Yӂ��F�	��*���l�l�%�y�w�}�W�������X��E�� ��l�%�y�u�w�}�Wϱ�����X��E�� ��l�:�6�1�{�}�W���Yӂ��GF�	��*���l�l�%�|�]�}�Wϸ�I����C9��Y��G���d�d� �g�m�>��������T��]�����3�8�
�g�$�n����&���F��Y��ʸ�%�}�u�u�w�}�>���G����F�N��;������h�w�q�W���Y����Z��`'��=��u�g�_�u�w�}�W���H����g.�	N�Y���u�u�u�1�"��>���Y���l�N�����4�u�_�u�w�}�W���I���G�� \�� ��e�
�e�_�w�}�W������F��G1�*���d�e�
�d�]�}�W���Y����W�	N����
� �d�e��-����s���F�S��U��!�%�b�
�"�l�G܁�K��ƓF�Q1�����
�g�&�f�9��(ށ�K����P	��X ��ʸ�g�e�f�������J���� T��h_�����u�0�0�<�w�<�W�ԜY���F��S�D�ߊu�u�u�u���#���Y���l�N��Uʱ�;�
���w�c�D��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��_�u�u�:�#�0����Y���F��^ �H���8�
�`�3��m�@���U���F�
��D��u�8�
�`�1��G���	��ƹF�N�����0�h�u�8��h����I�ѓ�C��RBךU���u�u�:�!�j�}����L����V��h�N�ߊu�u�
�
�4�-�Dݰ�&�Ԣ�lW��h;�U���:�%�;�;�w�m�3��M����l ��G1����g�&�d�d�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�t�W���	����^��d��U���u�1�;�u�i�)���&����W��G^�U���u�u�1�;�w�c����Nʹ��lW��1��Y���u�u�u�:�4�9�W�������
9��h_�D���6�1�y�u�w�}�WϺ������hY�����e�d�%�|�]�W�}���Y���G��T�����&�4�0�}�'��(���PӉ��G��D��ʸ�6�<�0�u�z�}�WϿ�&����@��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���%��
�&�w�`����-����l ��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�$�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���4�'������������9��R1�����a�l�4�&�0�}����
���l�N��������:�#�(�(��&ù��9��P1�L���&�2�
�'�4�g�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�4�
�>�����J����[��N��U���u�u�u�u�>�}�_���&�ғ�F9�� \��D��4�
�:�&��+�(���Y����l�N��U���u�u�u�u�w�<����<����x	��G��G���e�0�e�'�0�i�N��Y����u#��u/����� �
�d�
�"�;��������
P��=N��U���u�u�u�u�w�1��������T9��S1�A���!�0�u�u�w�}�W���Y���F���*������ �'�)�E���I����l��hZ�U��4�'������������9��Q��*���0�
�l�f�]�}�W���Y���F�R�����!�%�l�
�"�l�@݁�H����C9��Y�����g�|�!�0�w�}�W���Y���F�N��U���
�����(����K�ѓ�l��h��*��u�h�4�'���5�������G9�� 1�����
�
�0�
�n�e�}���Y���F�N�����3�}�!�%�n����N����[��G1�����9�g�d�|�#�8�W���Y���F�N��U���u�'�
����<���	����Q��h��*���
�c�u�h�6�/�1���;����F��C1�B���3�0�
�
�2��N��s���F�N��U���0�1�<�n�w�}�W���Y����]��QU��U���u�u�0�1�>�f�W�������A	��D����u�x�4�'���5�������G9�� 1�����'�2�a�g�6�.��������@H�d��Uʴ�'�����2����&����9��1����g�4�&�2��/���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u�6���������O��_��U���u�u�u�u�w�}����Q����
R��R	��L��h�4�
�:�$��݁�P�Ƹ�V�N��U���u�u�u�u�w�}����?����r%��B����b�e�0�d�%�:�C��E�ƭ�A9��r*��6���!� �
�d��(����K����lT��UךU���u�u�u�u�w�}����Yۇ��@��U
��@��u�=�;�_�w�}�W���Y���F�N��������:�#�(�(��&ù��9��P1�G��u�'�
����<���	����Q��B�����'�2�g�a�l�}�W���Y���F������}�8�
�a�%�:�E��Y�ƭ�l��D��؊�|�u�=�;�]�}�W���Y���F�N���������8�)����HĹ��V9��E��A��i�u�'�
���6�������lT��h�����a�'�2�g�a�f�W���Y���F�N�����u�}�8�
�c�/���@���R��X ��*���
�|�u�=�9�W�W���Y���F�N��Uʴ�'�����2����&����9��1����g�i�u�'���3���2����F��Y�� ���'�f�'�2�e�h�L���Y���F�N��U���u�3�_�u�w�}�W���Y����Z ��=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�'�
����<���	����Q��h^��*؊�0�
�e�u�$�4�Ϯ�����F�=N��U���
�����(����K�ѓ�lV��h\�����e�
�&�<�9�-����Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��-��������R�������u�u�u�u�w�}�WϷ�Yۇ��@��U
��G��|�!�0�u�w�}�W���Y���F�N���������"�-���N����lV��h��*��u�h�4�'���5�������G9�� 1�����l�'�2�a�a�W�W���Y���F�N�����}�%�&�2�5�9�E��PӒ��]FǻN��U���u�u�u�u�w�}����<����p-��C��*��
�
�
�
��8�(��Y����A��r+��4��� �%�!�g�`�8�G���J����U��h����u�u�u�u�w�}�W���Y����F�N��U���0�1�<�n�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����u#��u/����� �
�d�
���(݁�����F��D��U���6�&�{�x�]�}�W���&����q'��X�� ���d�
�
�
������@ù��@��h����%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �V�����1�
�d�`�w�5����Y���F�N��U���}�%�&�2�5�9�E��PӒ��]FǻN��U���u�u�u�u�w�}����<����p-��C��*��
�
�
�
��8�(��Y����A��r+��4��� �%�!�g�`�n����O����lR��d��U���u�u�u�u�w�8����Q����Z��S
��D��u�=�;�_�w�}�W���Y���F�N��������:�#�(�(��&����9��E��@��i�u�'�
���6�������lT��h��*ۊ�
� �d�c��n�}���Y���F�N�����<�n�u�u�w�}�W�������U]�N��U���0�1�<�n�w�}����	����@��=N��U���4�'������������9��1��G���2�`�e�4�$�:�W�������K��N���������8�)����HĹ��9��1�����e�4�&�2��/���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u�6���������S�C�����u�u�u�u�w�}�W���Q����Z��S
��D��u�=�;�_�w�}�W���Y���F�N��������:�#�(�(��&����9��E��@��i�u�'�
���6�������lT��h��*؊�0�
�g�n�w�}�W���Y���F��[��U´�
�<�
�1��l�A������F�N��U���u�u�u�u�6�/�1���;����F��C1�B���e�g�g�'�0�h�G��Y����u#��u/����� �
�d�
���(܁�����9��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�3�u�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�����w$��|�����g�b�0�e�d�o����L����@��YN�����&�u�x�u�w�<����<����x	��G��G���0�e�f�g�%�:�B�������]9��X��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ����D�����g�a�|�!�2�W�W���Y���F�N��U´�
�<�
�1��l�O������F�N��U���u�u�u�u�6�/�1���;����F��C1�B���e�f�g�'�0�h�G��Y����u#��u/����� �
�d�
���(���&����9F�N��U���u�u�u�9�>�}��������W9��X�����u�u�u�u�w�}�W���Y�����h(��1���� �%�!�e�j����J�ԓ�V�� ^��Hʴ�'�����2����&����V9��1�����f�m�%�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C���������"�-���N����lV��h��*��u�&�<�;�'�2����Y��ƹF��E��0����� �%�#�o�@���H�֓�l��h[�*���<�;�%�:�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�%�&�0�?���M����[��N��U���u�u�u�u�>�}��������W9��V�����u�u�u�u�w�}�W���Y�����h(��1���� �%�!�e�j����I�ԓ�V��^��Hʴ�'�����2����&���� 9��1�����f�m�_�u�w�}�W���Y���V
��QN�����2�7�1�g�c�t����Y���F�N��U���u�u�u�'���3���2����F��Y��*ۊ�
�
�0�
�a�}�JϿ�����w$��|�����g�b�0�d�g�n����M�ޓ� ]ǻN��U���u�u�u�u�9�}��ԜY���F�N��ʼ�n�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����<����p-��C��*��
�
�
�
��8�(��Y����T��E�����x�_�u�u�%��2���8����G��h\�*���
�
�
�0��h�(�������A	��N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W����έ�l��h��*��`�u�=�;�w�}�W���Y���F��QN�����2�7�1�g�c�t����Y���F�N��U���u�u�u�'���3���2����F��Y��*ۊ�
�
�0�
�b�}�JϿ�����w$��|�����g�b�f�0�f�k����J����F�N��U���u�u�0�&�1�u��������lT��G�����_�u�u�u�w�}�W���Y���R��q+��7���:�!� �
�f��(ށ�&����T9��N�U���
�����(����K�ѓ�lW��h]�� ��a�
�f�_�w�}�W���Y���F��SN��N���u�u�u�u�w�8�Ϸ�B���F�N��ʼ�n�u�u�0�3�-����
��ƹF�N��������:�#�(�(��&����9��E��@��4�&�2�u�%�>���T���F��E1��0����:�!� ��l�(���&����A��Z�����2�
�'�6�m�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�4�
�<��9�(��L�Ƹ�VǻN��U���u�u�u�u�1�u��������lT��G�����_�u�u�u�w�}�W���Y���R��q+��7���:�!� �
�f��(ށ�&����T9��N�U���
�����(����K�ѓ�lW��h��*��n�u�u�u�w�}�W���YӃ��Z �V�����1�
�d�c�w�5��ԜY���F�N��U���u�4�'����4�������W��R1��G���'�2�`�e�k�}����<����p-��C��*��
�
�
�
��(�F��&����F�N��U���u�u�0�1�>�f�W���Y���F��Y
�����u�u�u�u�2�9���Y����]��E����_�u�u�x�6�/�1���;����F��C1�B���d�f�g�'�0�h�GϿ�
����C��R��U���u�u�4�'���5�������G9�� 1��D���g�'�2�`�g�<����&����\��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}��������T9��S1�A���!�0�_�u�w�}�W���Y���Z �V�����1�
�d�m�w�5��ԜY���F�N��U���u�4�'����4�������W��R1��F���'�2�`�e�k�}����<����p-��C��*��
�
�
�
�2��A��Y���F�N��U���9�<�u�4��4�(���&����F��R ��U���u�u�u�u�w�}�W�������v#��v-�� ���!�g�b�0�f�n�E�������Z�V��3�����:�!�"��F؁�&¹�� 9��h_�E���n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�;�w�;�W���Y����������u�;�u�'�4�.�L�ԜY�����h �����'�
�d�
��8�(��Y����T��E�����x�_�u�u�%���������W��^1�����l�4�&�2��/���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F��QN�����2�7�1�c�`�}����s���F�N��U���u�u�4�'�9�9�(�������l��R	��D���h�4�
�:�$��݁�B���F�N��U���u�9�<�u�6���������W�C��U���u�u�u�u�w�}�W���YӇ��l��R1�����d�
�
�0��l�W������\��C��*��
�
�
� �f�i�(��s���F�N��U���0�1�<�n�w�}�W���Y����]��QU��U���u�u�0�1�>�f�W�������A	��D����u�x�6�
���6�������V��h^�����e�u�&�<�9�-����
���9F���<�����!�'��o�(���&����V��V�����'�6�o�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�WϷ�Yۇ��@��U
��@��u�=�;�_�w�}�W���Y���F�N��*������0�:�o�G���I����lQ��R���������8�)����HĹ��9��1����e�_�u�u�w�}�W���Y�Ʃ�@�������7�1�g�`�~�)����Y���F�N��U���u�u�9����%�������9��1����`�i�u�'���3���2����F��Y��*���
�
�0�
�c�f�W���Y���F�N�����3�_�u�u�w�}�W����ƥ�FǻN��U���;�u�3�_�w�}��������@]ǑN��X���9�����)����Kù��9��P1�Bʴ�&�2�u�'�4�.�Y��s���P
��y*��4���0�8�g�e�2�l����O�ѓ�@��Y1�����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�;�_���
����W�� _�����u�u�u�u�w�}�W���Y�����~ ��-���!�'�
�g���(���&����[��E��0����� �%�#�o�@���H�֓�l��h[�N���u�u�u�u�w�}�Wϻ�
���R��^	�����d�`�u�=�9�W�W���Y���F�N��Uʶ�
�����8���I����l��hX�U��4�'������������9��R1��L���2�f�m�_�w�}�W���Y���F��SN��N���u�u�u�u�w�8�Ϸ�B���F�N��ʼ�n�u�u�0�3�-����
��ƹF�N��*������0�:�o�E���I����lP�������%�:�0�&�w�p�W�������w#��e<�����g�
�
�
�2��N܁�
����l��TN����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�<�u�6���������O��_�����u�u�u�u�w�}�W���Y����}"��v<�����g�g�0�e�%�:�A��E�ƭ�A9��r*��6���!� �
�d���(ށ�&����_��=N��U���u�u�u�u�w�1��������T9��S1�@���!�0�u�u�w�}�W���Y���F���<�����!�'��o�(���&����_��S���������"�-���N�Փ�lV��h��*��n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�;�w�;�W���Y����������u�;�u�'�4�.�L�ԜY�����~ ��-���!�'�
�g���(���&����R��P �����&�{�x�_�w�}����=����a��Z1�G���d�'�2�c�b�<����&����\��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���3�}�%�&�0�?���H�Ƹ�V�N��U���u�u�u�u�w�}����7����a4��E��G؊�
�
�0�
�c�}�JϿ�����w$��|�����g�b�0�d�f�o����L����F�N��U���u�u�0�&�1�u��������lT��G�����_�u�u�u�w�}�W���Y���P
��y*��4���0�8�g�g�2�l����O���F��E1��0����:�!� ��l�(܁�&¹��A��V����u�u�u�u�w�}�W���Y����F�N��U���0�1�<�n�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����}"��v<�����g�a�0�e�%�:�A������]F��X�����x�u�u�6���2���+����lT��h��*���
�m�
�&�>�3����Y�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��U´�
�<�
�1��j�^Ϫ���ƹF�N��U���u�u�u�u�;��3���+����^9��1��E���2�c�d�i�w�/�(���=����\��B��D݊�
�
�
�
�2��O��Y���F�N��U���9�<�u�4��4�(���&����F��R ��U���u�u�u�u�w�}�W�������w#��e<�����g�
�
�
�2��O���DӇ��l ��s,��>���%�!�g�b�2�m�E�������l�N��U���u�u�u�0�3�4�L���Y���F���U���u�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�>�(���<����G��h\�*���
�0�
�f�w�.����	����@�CךU���9�����)����Kǹ��9��P1�F���&�2�
�'�4�g�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y����UF��G1�����1�`�d�u�?�3�}���Y���F�N��U���6�
��������K�ғ�lW��R	��F���h�4�'����4�������W��R1��G���'�2�`�e�]�}�W���Y���F�R�����%�&�2�7�3�o�B�������9F�N��U���u�u�u�u�w�1�>���!����V��\�����'�2�c�f�k�}����<����p-��C��*��
�
�
�
�2��@��Y���F�N��U���;�u�3�_�w�}�W���Y�Ʃ�WF��NךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�9����%�������9��1����l�4�&�2�w�/����W���F�T��;�����0�8�e�k��������_��D�����:�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Q����Z��S
��B���!�0�u�u�w�}�W���Y���F���<�����!�'��o�(���&����P��S���������"�-���N����lU��h��*��n�u�u�u�w�}�W���YӃ��Z �V�����1�
�d�`�w�5��ԜY���F�N��U���u�6�
����%�������l��h��*��u�h�4�'���5�������G9�� 1��E���'�2�a�e�]�}�W���Y���F�R ����u�u�u�u�w�}�������F�N�����<�n�u�u�2�9��������9F�C��������2�0�E����ד�V��_�����;�%�:�0�$�}�Z���YӅ��z(��o/�����
�g�
�
��8�(��&����T��E��Oʥ�:�0�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��|�!�0�_�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�<�w�<�(���&����Q�����ߊu�u�u�u�w�}�W���Y�Ư�l/��r6��'���8�g�c�0�f�/���H���R��q+��7���:�!� �
�f��(ށ�&����T9��UךU���u�u�u�u�w�}����Yۇ��@��U
��G���|�!�0�u�w�}�W���Y���F�N��������!�%��Eف�&¹��T9��N�U���
�����(����K�ѓ�lW��h��*��n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�;�w�;�W���Y����������u�;�u�'�4�.�L�ԜY�����E��C��4�&�2�u�%�>���T���F��h��*��
�&�<�;�'�2�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}�'�.��������O��_��U���u�u�u�u�w�}��������T9��S1�A���!�0�u�u�w�}�W���Y���F������c�e�i�u�'�>�����Փ�l�N��U���u�u�u�0�$�;�_���
����W��Z�U���;�_�u�u�w�}�W���Y���F��h��*��u�h�<�g�1��E���	��ƹF�N��U���u�u�;�u�1�W�W���Y���F��SN��N�ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�e�/���AӇ��Z��G�����u�x�u�u�>�����O˹��@��h����%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�>�}��������W9��_�����u�u�u�u�w�}�W���Y�����E��L��i�u�%�6�9�)����I���F�N��U���u�0�&�3��-��������S�����ߊu�u�u�u�w�}�W���Y�ƥ�l��hW�U��<�f�3�
�b�d���Y���F�N��U���;�u�3�_�w�}�W���Y�Ʃ�WF��NךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�f�'�0�d�NϿ�
����C��R��U���u�u�<�
�2��@ց�
����l��TN����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�<�u�6���������S�C��U���u�u�u�u�w�}�W���Yӏ��A��Y�I���%�6�;�!�;�o�G�ԜY���F�N��Uʰ�&�3�}�%�$�:����K������YNךU���u�u�u�u�w�}�W���J����l_��R�����3�
�c�l�'�f�W���Y���F�N�����3�_�u�u�w�}�W����ƥ�FǻN��U���;�u�3�_�w�}��������@]ǑN��X����9�
�:��2��������Q��D��ʥ�:�0�&�u�z�}�WϷ�&����\��X�����2�l�b�4�$�:�(�������A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�o�^������F�N��U���u�u�u�u�>���������C9��E��L��i�u��9��2�(���	����A��_�N���u�u�u�u�w�}�Wϻ�
���R��^	�����d�b�u�=�9�W�W���Y���F�N��Uʼ�
�<��'��2�(�������F������!�9�f�e�]�}�W���Y���F�R ����u�u�u�u�w�}�������F�N�����<�n�u�u�2�9��������9F�C����2�a�m�4�$�:�W�������K��N�����2�a�m�4�$�:�(�������A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��U���u�u�u�<�%�:�C��E�ƥ�9��P1�M��u�u�u�u�w�}�W�������N��h��*���
�f�|�!�2�}�W���Y���F�N��U���
�0�
�`�w�`��������_��UךU���u�u�u�u�w�}�������F�N��Uʰ�1�<�n�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z���
������T��[���_�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�3�8�g�~�}����Y���F�N��U���'�
������������lU��h^��D���2�f�a�u�j�<����<����x	��G��G���f�0�e�d��(�F��&����F�N��U���u�u�4�'���5�������G9�� 1�����g�'�2�f�e�}�JϿ�����w$��|�����g�b�f�0�g�o����H�ӓ� ]ǻN��U���u�u�u�u�%��2���8����G��h\�*ي�
�
�
�0��m�C��Y����u#��u/����� �
�d�
���(ځ�����
9��d��U���u�u�u�u�w�<����<����x	��G��G���f�0�e�m�%�:�D��Y����A��r+��4��� �%�!�g�`�n����A����W��h����u�u�u�u�w�}�W���&����l��h]�A��u�0�
�8�e�;�(��N����9F�N��U���u�u�u�0��0�C�������F���*���a�3�
�d�g�-�L���Y���F�N��U���
�8�
�0��m�O��Y����G��Q��E���%�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���Ĺ��^9����U´�
�:�&�
�!��W�������]��Q��A���%�|�|�!�2�W�W���Y���F�N��������:�#�(�(��&����9��h��*��e�i�u�'���3���2����F��Y��*���
�`�3�
�b�k���Y���F�N��U���'�
������������lU��h_��@���2�f�d�u�j�<����<����x	��G��G���f�0�d�d��(�F��&����F�N��U���u�u�6�
�#���������l��h��*��`�i�u�9�;���������9��1��*���d�%�n�u�w�}�W���Y�����[�����:�%�g�
������K���F��h��3����:�
�`�2�l����L�ד� ]ǻN��U���u�u�u�u�;�1�(���&����lT��R1�����f�g�u�h�4���������C9��h��*���d�l�
�f�]�}�W���Y���F�T�����'��:�
�`�8�F�������F������:�
�:�%�e��(ށ�����9��d��U���u�u�u�u�w�>�(���?����\	��[��*ڊ�0�
�g�c�k�}����&����	��h]�����3�
�c�f�'�f�W���Y���F�N�����
�:�
�:�'�n�(���&���� T��R�����!��'��8��B���H����P��h����u�u�u�u�w�}�W�������A9��X��D���2�f�a�u�j�;�(���?����\	��_�� ��f�
�f�_�w�}�W���Y���F��h��3����:�
�f�%�:�D��Y����`9��h(��*���%�f�
� �f�h�(��s���F�N��U���&�9�!�%�a�/���M�����h��D܊� �d�b�
�e�W�W���Y���F�N�����%�b�'�2�d�k�W��
����^��h��D��
�g�_�u�w�}�W���Y���@��C��M���2�f�b�u�j�.����	�ޓ�F9��^��G�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�C������F��R ךU���u�u�u�u�w�}����<����p-��C��*��
�
�
�
��8�(��Y����A��r+��4��� �%�!�g�`�n����A����lU��UךU���u�u�u�u�w�}����<����p-��C��*��
�
�
�
��8�(��Y����A��r+��4��� �%�!�g�`�n����H¹��T9��Z�U���u�u�u�u�w�}����?����r%��B����b�f�0�d�a�/���O���R��q+��7���:�!� �
�f��(���&˹��lW��1��N���u�u�u�u�w�}�WϿ�����w$��|�����g�b�f�0�f�d����J���F��E1��0����:�!� ��l�(܁�&¹��l ��\�*��_�u�u�u�w�}�W���Y����u#��u/����� �
�d�
���(���&����[��E��0����� �%�#�o�@����֓�l��h]�A�ߊu�u�u�u�w�}�W�������v"��t%�����
�d�
�
������H�����h(��1���� �%�!�e�j�D���I�ԓ�V��\����u�u�u�u�w�}�W���&����q'��X�� ���d�
�
�
��8�(��Y����A��r+��4��� �%�!�g�`�n����L����T��h����u�u�u�u�w�}�W���&����q'��X�� ���d�
�
�
��8�(��Y����A��r+��4��� �%�!�g�`�n����K����W��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���R�������!�9�d�e�j�8�����ד�F9��]��G���;�u�4�
�8�.�(���&���G��^�����`�`�%�|�~�)��ԜY���F�N��Uʴ�'�����2����&����Q��R��U��4�'�9�
�8�����JŹ��V9��Z�� ��d�
�f�_�w�}�W���Y���F��E1��0����:�!� ��l�(�������Z�V�����:�
�:�%�d��(���&�ғ�F9��_��F�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�l�JϿ�&���R��Y��]���&�4�!�h�6�����&����P9��G�����_�u�u�u�w�}�W���Y����u#��u/����� �
�d�
�"�;��������
R��S���������"�-���N����U�� UךU���u�u�u�u�w�}����<����p-��C��*��
� �3�'�e�/���L�����h(��1���� �%�!�e�j��������9F�N��U���u�u�u�'���3���2����F��Y�� ���'�f�'�2�e�h�W������v#��v-�� ���!�g�b�7�1�8�(��Y���F�N��U���'�
������������l��Q��A���2�g�c�u�j�<����<����x	��G��G���7�3�0�
�l�}�W���Y���F���*������ �'�)�E�������A9��E��G��u�h�4�'���5�������G9�� 1�����
�n�u�u�w�}�W���Y����A��r+��4��� �%�!�g�`�?����&Ź��T9�� ]��Hʴ�'�����2����&����Q��R��N���u�u�u�u�w�}�WϿ�����w$��|�����g�b�7�3�2��(���&����Z�V��3�����:�!�"��F؁�����lT��N��U���u�u�u�u�6�/�1���;����F��C1�B���3�0�
�
�2��N��E�ƭ�A9��r*��6���!� �
�d��(����J���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���f�3�8�g�~�<����	����@��A_��U���-�!�:�1��(�E��&���R�������!�9�g�g�j�)���J����S��h�\���=�;�u�u�w�}�W���Y����A��r+��4��� �%�!�g�`�?����&�����h��3����:�
�c�d�8�G��&����W��G]�U���u�u�u�u�w�}����?����r%��B����b�7�3�0��}�JϿ�����u	��{��*���f�0�d�d��(�E��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�f�3�8�e�t����Q����\��h��*���u�-�!�:�3����O����F��SN�����%�6�;�!�;�o�E������U��B1�Bߊ�d�|�4�1�9�)�_�������l
��h_��U���
�e�
� �e�j�(��PӇ����F��*���&�
�#�
�w�}����I����lT��1��\���u�=�;�u�w�}�W���Y�����h(��1���� �%�!�e�j��������[��E�����'��:�
�a�n����Hǹ��lT��1��N���u�u�u�u�w�}�WϿ�����w$��|�����g�b�7�3�2��W������G9��E1�����c�f�0�d�f����O¹��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�f�3�:�o�^Ͽ��έ�l��D��ۊ�u�u�-�!�8�9�(���K����CT�V ��]���6�;�!�9�e�m�JϪ�	����l ��[�*��|�u�=�;�w�}�W���Y���F��E��0����� �%�#�o�@�������F���*����'��:��k�D���H����U��X����u�u�u�u�w�}�W�������v#��v-�� ���!�g�b�7�1�8�(���DӇ��l
��q��9���
�c�f�0�g�l�(���K����CU��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�a�1�0�E������R��X ��*���
�u�u�-�#�2����&����l����U´�
�:�&�
�!��W�������9��h\�@���|�|�!�0�]�}�W���Y���F�V��3�����:�!�"��B��E�ƭ�A9��S�����m�
�:�1�'�4����N�ߓ� ]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�W���Y������C��ߊ� �d�c�
�e�`��������_��G��\ʡ�0�_�u�u�w�}�W���Y�ƭ�A9��r*��6���!� �
�`�g�1��������
^�
N��������:�#�(�(���I���F�N��U���u�4�'����4�������S��h�����2�f�e�u�j�<����<����x	��G��Mߊ�n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���M����lT����U´�
�:�&�
�!��W�������]��B1�Lي�g�u�;�u�8�u��������_��N�����d�a�3�
�`�h����P�Ƹ�VǻN��U���u�u�u�u�%��2���8����G��hV��D��u�'�
�:�2�)����H����W9��^1��*��l�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���=�;�u�u�w�}�W���Y����A��C1�����:�
�m�f�2�m�F߁�����W�
N�����
�:�
�:�'�o�(܁�&ù��l ��W�*��_�u�u�u�w�}�W���Y����_��X�����g�
�
�
������K���F��E1��*���
�:�%�g���(߁�&����
V��G]�U���u�u�u�u�w�}��������A9��X��M���0�e�a�'�0�n�N���DӇ��l
��q��9���
�m�f�0�g�i����@�ғ� ]ǻN��U���u�u�u�u�%���������C9��h]��*ڊ�
�0�
�g�a�a�W���&����\��X��GҊ�
�
�
�
�"�l�Dځ�J���F�N��U���u�4�'�9��2�(���	���� 9��1�*���
�f�d�i�w�/�(���?����\	��V��*���
�e�3�
�g�d���Y���F�N��U���'�
�!��%�����A�Փ�lW��h��*��c�i�u�'��)�1���5����^��h��*ۊ� �d�c�
�d�W�W���Y���F�N�����
�:�
�:�'�o�(܁�&¹��A��]�U��4�'�9�
�8�����K˹��V9��1��*��b�%�n�u�w�}�W���Y�����h��3����:�
�m�d�8�F������� W��S�����!��'��8��O����ד�l ��W�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����W�N���ߊu�u�u�u�w�}�W�������l ��h"����
�
�
�
��8�(��Y����A��C1�����:�
�c�f�2�m�C���&����l��=N��U���u�u�u�u�w�/�(���?����\	��X��*���
�0�
�c�w�`��������A9��X��C���0�e�d�3��i�F���B���F�N��U���u�'�
�!��/�;���&�Г�l��h\�����g�u�h�4�%�1�(���&����lU��1��D���3�
�`�c�'�f�W���Y���F�N�����!��'��8��A����ד�V��W��Hʴ�'�9�
�:��2���&����9��Q��@���%�n�u�u�w�}�W���Y����A��C1�����:�
�c�0�g�o��������Z�V�����:�
�:�%�d��(���&Ĺ��lT��1��N���u�u�u�u�w�}�WϿ�����u	��{��*���0�e�f�&�%�:�O��E�ƭ�A9��h(��*���%�f�
�
���F���&����l��=N��U���u�u�u�u�w�/�(���?����\	��X��*ۊ�
�
�0�
�d�}�JϿ�����u	��{��*���f�0�d�b�1��B���	��ƹF�N��U���u�u�'�
�#���������l��h]��*���
�a�u�h�6�/��������\��1�����d�
� �g�b��D�ԜY���F�N��Uʴ�'�;�1�
�2�0�Oށ�&����T��S�����!��'��8��E���M����U��h����u�u�u�u�w�}�W���&����l��Z1�*ۊ�0�
�d�u�j�<����&����	��h\��F���3�
�f�m�'�f�W���Y���F�N�������!�'��k�(���&����P��S�����!��'��8��O����֓�l��h]�C�ߊu�u�u�u�w�}�W�������w*��R��D���0�d�'�2�o�n�K�������l ��h"����
�
�
�
��8�(��O���F�N��U���u�6�
� ������H�ߓ�lT��R	��B���h�4�'�9��2�(���	���� 9��1�����f�l�n�u�w�}�W���Y�����u;��9���'�
�c�
������K�����h��3����:�
�m�d�8�F������� W��=N��U���u�u�u�u�w�1�5���5����^9��1��A���2�b�l�i�w�/�(���?����\	��V��*���
�
�0�
�e�k�}���Y���F�N����� ���0�:�l�N���L����l^��R�����9�
�:�
�8�-�Eׁ�&����9��P1�D��u�u�u�u�w�}�W�������}"��C��*��
�
�
�0��m�W������G9��E1�����m�f�0�e�f�����J����F�N��U���u�u�6�
���2�������l��h��*��u�h�4�'�;���������9��R1��Dڊ�0�
�f�d�]�}�W���Y���F�T�� ����0�8�d�n�8�G�������Z�V�����:�
�:�%�e��(؁����� 9��d��U���u�u�u�u�w�>�(���=����A�� W��*ۊ�0�
�`�u�j�<����&����	��h\��F��
� �g�f��n�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�6�.��������@H�d��Uʥ�:�0�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��|�!�0�_�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C[�����|�4�1�}�'�>�����ד�[��O�����
� �d�f��o�^�����ƹF�N��U���u�u�'�
�8�8����&����9��E��@��i�u�'�
�8�8����&���� 9��Q��G���%�n�u�u�w�}�W���Y����A��X
�����
�d�
�
��8�(��Y����A��X
�����
�d�
�
��(�F��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�f�t�^Ϫ����F�N��U���u�3�
���	����O����lU��N�U�������#�h�(���K����CU��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�f�1�0�F���PӒ��]l�N��U���u�u�u�3���;���6����9��E��F��u�h�3�
���E�������9��h_�D���n�u�u�u�w�}�W���YӒ��lP��E��F��u�h�!�%�a����@ǹ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�e�3�:�d�^�����ƹF�N��U���u�u��-��$����L����lU��N�U���
� �l�d�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9�� 1����|�u�=�;�w�}�W���Y���F��{1��*���
�:�%�d��8�(��A���Z*��^1�����:�
�c�3��i�E���B���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������A	��D�X�ߊu�u�'�6�$�}������ƹF��R	�����u�u�u�3��-���������������h�r�r�u�?�3�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�d�|�w�5����Y���F�N��U���
�0�
�l�a�a�W���&����P��G\�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��B���8�d�|�|�w�5����Y���F�N��U���
�e�b�i�w�/�(���@�ד�]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�b�1�0�F���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�|�!�0�]�}�W���Y���F�E��D��u�h�2�%�1��Nځ�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���d�3�8�g�~�t����s���F�N��U���&�9�!�%�f�4����J����[��R����
�
� �g�d��E�ԜY���F�N��Uʦ�9�!�%�e�>�/���L�����h��Gڊ�
� �g�c��o�}���Y���F�N�����!�%�l�<�%�:�D��Y����V
��Z�*��� �g�m�
�e�W�W���Y���F�N�����%�b�<�'�0�n�A���Dӕ��l��Y��*���g�m�
�g�]�}�W���Y���F�C��Bފ�0�
�f�b�k�}����M����T��h����u�u�u�u�w�}�W���&�֓�V��Z�I���8�
�e�3��o�@���B���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������A	��D�X�ߊu�u�'�6�$�}������ƹF��R	�����u�u�u�3��-���������������h�r�r�u�?�3�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�d�u�9�}��������l ��^�*��h�4�
�:�$��ށ�P����[��N��U���u�u�u�u�#�-�Nہ�����
W�
N����
� �d�b��l�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�#�8����Y����VF��G1��*���|�:�u�=�w�)��������VH�d��Uʴ�
��3�8�6�.���������T��U´�
�!�'�y�6��$����ƭ�l�������!�e�'�4��8����&����CT�R�����`�3�
�e�g�-�[ϻ�����WR��B1�Fފ�g�u�-�!�8�9�(���H����CT�R�����g�3�
�a�a�-�[ϻ�����WW��B1�Cي�g�u�-�!�8�9����O�Փ�OǻN�����_�u�u�u�w�<�Ͽ�&����@��Dd��U���u�u�u�"�2�}����&����U��N��U���u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y������D����4�
�:�&��2����P���G��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d�1�0�G�ԜY���F�N��Uʰ�1�<�n�u�w�}�W���Yӑ��]F��h=�����3�8�d�h�w�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�-�!�:�3����Où��[��G1�����9�d�e�|�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��A�ߊu�u�u�u�w�}�W�������N��G1�����9�2�6�d�j�<�(���Y������C��ߊ� �d�c�
�e�`��������_��G��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�n����K���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!��.�(���G���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�u�u�0�$�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}�������F�N��Uʢ�0�u�%���)�(���&���l�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
�ԓ�@��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��F�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���&����F�d��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Qۇ��P	��C1��D��h�0�<�6�9�i����K�ғ�O�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!��.�(��Y���F�N��U���9�<�u�}�6�����&����P9��
N��*���u�;�u�4��2����¹��F��^�����3�
�g�a�'�t�^Ϫ����F�N��U���u�u�u�4������E�ƭ�l5��D�����a�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��h��*���k�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��Y1�����e�'�4�
�2�9����H����[��G1�����9�d�e�u�%�3����	����@��A_��U���-�!�:�1��(�F��&���O�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}�>�����&ù��R��R�����d�
�g�h�6�����&����O�V ��]���6�;�!�9�f�m�Jϻ�����WU��B1�BҊ�g�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
�Г�@��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��@�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���&����F�d��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Qۇ��P	��C1��D��h�0�<�6�9�o����M�Г�O�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�d�;���B���F�N��U���u�9�<�u��<�(���
����T��N�����0�u�;�u�6�����&����F�R�����g�3�
�a�a�-�^�������F�N��U���u�u�u�u�6��$������R��c1��M���8�b�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӈ��`2��CV�����u�k�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����*����Z�V��!���l�3�8�m�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��ӊ�&�
�u�k�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������l ��R������&�d�
�$��L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�d����A���F�N��U���u�0�1�<�l�}�W���Y�����YN��*���&�d�
�&��}�I�ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$����֓�@��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���;�4�
��$�l�(���&���FǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����l ��h_����u�u�u�u�w�}�W������F�N��U���u�u�u�%������DӇ��`2��C_�����d�n�u�u�w�}�W���Y����]��QUךU���u�u�u�u�?�3����-����9��Z1�U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��Dي�&�
�g�_�w�}�W���Y���F��DךU���u�u�u�u�w�}�W���	����U��S�����
�!�g�3�:�l�L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:�����3�8�d�u�i�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d��.�(��s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!�c�;���Y���F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���Hƹ��^9��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$����ӓ�@��N��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�%������DӇ��`2��C_�����d�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�c�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�`�h�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�b�3�:�l�L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���u�u�0�1�>�f�W���Y���F��_������&�d�
�$��A��Y���F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	���&����Q�	NךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�d�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��1����u�k�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����*����Z�V��!���g�
�&�
�n�W�W���Y���F�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�n�;���B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�e�3�8�f�}�I�ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�o�(���&����F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$����֓�@��UךU���u�u�u�u�w�}�������F�N��Uʢ�0�u�%���)�F�������X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�
���F�N��U���u�u�u�4������E�ƭ�l5��D�*���
�e�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����T��D��D��u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��݊�&�
�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�g�
�&��l�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��Gي�&�
�g�h�w�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�f�m�Jϻ�����WW��B1�Cي�g�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��\�U���u�u�u�u�w�}�������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��h�����#�
�u�u�/�)����&����P��G\��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Eہ�
����l�N��U���u�u�u�0�$�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����l ��h\����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���������� F�d��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Qۇ��P	��C1��D��h�0�<�6�9����@����O������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d�1�0�G�ԜY���F�N��Uʰ�&�3�}�}�'�>��������lW������4�1�}�%�4�3����H�����C�����
�c�f�%�~�t����s���F�N��U���u�u�4�
��;���Y����g9��Z�����f�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���a�3�8�g�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӊ��V��
P�����u�u�u�u�w�}�W���7����^F�L��-���������/���!����F�N�����6�&�n�u�w�8�Ϯ�����lǻN��Xʴ�
�:�0�4�$�:�W�������K��N�����:�0�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^����0�u�%�&�0�>����-����9��Z1�Yʰ�<�6�;�
�"�o�N܁�K���F��P��U���u�u�<�u��3����	����@��X	��*���u�%�&�4�#�t����Q����\��h�����u�u�%�&�0�>����-����l ��h^��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�a�3�:�o�^Ͽ�ӈ��N��h�����#�
�u�u�/�)��������
U��G��\���=�;�_�u�w�}�W���Y����\��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��2���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������@��YN�����&�u�x�u�w�<�(�������Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�~�}�Wϼ���ƹF�N�����;�!�}�%�4�3��������[��G1�����|�4�1�}�'�>��������lW������6�0�
��$�l����I���G��d��U���u�u�u�4��9���Y����\��h�����n�u�u�u�w�8����Y���F�N�����9�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�'�4�.�<����Y����V��C�U���4�
�0�1��.����	����	F��X��´�
�0�u�%�$�:����&����GT��Q��G���0�<�6�;��(�E��&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���������� O��Y
�����4�
�:�&��+�(���Y����P	��h��G��
�g�|�|�#�8�W���Y���F������,�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������R��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�ƭ�l��B��E��u�9����)����Oʹ��9��P1�@�ߊu�u�%�'�#�/�(���DӅ��q3��{+�����c�
�
�
�2��F��Y����C9��C��*���h�6�
� ������H�ߓ�lT��R	��B��u�u�4�
�2�(���E�Ư�l$��s"�����d�l�0�f�%�:�O��s���R��R����i�u�9�������&����V9��E��B��_�u�u�%�%�)����Y����_9��y*�����
�c�
�
��8�(��B�����E�����u�h�6�
���2�������l��h��*��n�u�u�4��8����N���P
��b ��0���8�d�l�0�`�/���@���F��h�� ���m�i�u�9���;�������
9��1����d�_�u�u�'�/����&�����u;��9���'�
�b�
������L��ƓF�C�����2�7�1�d�o�<����Y����V��C�U���4�
�<�
�3��Gׁ�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&����T��X����|�n�u�u�2�9��������9l�N�U���&�2�7�1�f�j�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����W��S�����:�&�
�#��}�W���:����^N��
�����d�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�l�OϿ�
����C��R��U���u�u�4�
�>�����K˹��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��]�����:�d�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�F������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�}���Y����]l�N��U���u�u�u�4��4�(���&����[������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�2�_ǿ�&����GF�V�����
�:�<�
�~�t�}���Y����C��R���ߊu�u�x�4��4�(���&������^	�����0�&�u�x�w�}��������W9��Y�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����b�b�i�u�6�����&����F�V��&���8�m�1�"�#�}�^��Y����]��E����_�u�u�x�w�-��������P��V�����'�6�&�{�z�W�W���	����l��h_�B���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�c�u�j�u��������EW��S�����
�&�}�d�3�*����H����F�R �����0�&�_�_�w�}�ZϿ�&����Q��Y�U���<�;�%�:�2�.�W��Y����C9��P1����b�
�&�<�9�-����Y����V��V��&���8�_�u�u�2�4�}���Y���F�N�����<�
�1�
�`�j�K�������]��[��D��4�
��3�:�l�W������O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��b�4�&�2�w�/����W���F�V�����1�
�b�b�6�.���������T��]����
�&�|�w�}�������F�N��U���u�%�&�2�5�9�F��Y���R��X ��*���
�u�u�%������Aӂ��]��V��N���u�0�1�%�8�8��Զs���K��G1�����1�g�a�u�$�4�Ϯ�����F�=N��U���&�2�7�1�e�i�(�������A	��N�����&�!�%�l��(�F��&���F�U�����u�u�u�u�w�}�WϿ�&����Q��_�U��}�:�}�!�'�d�(���H����CW������!�9�g�g�~�<�ϰ��θ�C9��h��D��
�d�h�4��2��������F��SN�����8�
�a�3��m�E���Y�ƭ�l��D��؊�|�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��l�BϿ�
����C��R��U���u�u�4�
�>�����H�ӓ�@��Y1�����u�'�6�&��-�������@��1�����0�1�3�
�f��E�ԜY�Ʈ�T��N��U���u�u�u�u�6���������S�
N�����:�&�
�:�>��W���	������ ��]¼�
�0�0�
��8��������lT��h�Hʴ�
�:�&�
�!��^���s���V��G�����_�_�u�u�z�<�(���&����W�������%�:�0�&�w�p�W�������T9��S1�A܊�&�<�;�%�8�}�W�������R��^	������
�!�
�$��[ϻ�����WU��B1�BҊ�g�_�u�u�2�4�}���Y���F�N�����<�
�1�
�f�k�K���Q����\��h�����u�u�%�&�0�>����-����l ��h[�����}�%�6�;�#�1�F��DӃ��G��S]�� ��b�
�g�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��AӇ��Z��G�����u�x�u�u�6���������^��D�����:�u�u�'�4�.�_���
����@��d:��ߊ�&�
�y�0�>�>�������� R��GךU���0�<�_�u�w�}�W���Y���R��^	�����d�m�i�u��-��������Z��S�����2�6�0�
��.�B������R��Y��]���6�;�!�9�f�m�Jϻ�����WR��B1�Fފ�g�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�o�B���
������T��[���_�u�u�%�$�:����K����R��P �����o�%�:�0�$�<�(���&����l5��D�����a�u�-�!�8�9�(���H����CT�N�����;�u�u�u�w�}�W���YӇ��@��U
��G���u�h�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����#�
�u�u�/�)����&����U��G\��N���u�0�1�%�8�8��Զs���K��G1�����1�g�`�u�$�4�Ϯ�����F�=N��U���&�2�7�1�e�h�(�������A	��N�����&�<�
�0�2��(�������W9��h\�*��u�%�&�2�4�8�(���
�ӓ�@��N�����;�a�3�
�e�i����Y����V��=N��U���u�u�u�u�w�-��������S��S��]���6�;�!�9�0�>�F������T9��R��!���`�3�8�a�w�3�WǷ�&����G9��E��*���1�3�
�d��o�JϿ�&����G9��1�U���u�:�}�4��2����¹��F��^�����3�
�g�a�'�t�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������_��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��_�*���<�;�%�:�w�}����
�έ�l��h�����
�!�f�3�:�o�[ϻ�����WW��B1�Cي�g�_�u�u�2�4�}���Y���F�N�����<�
�1�
�f�d�K���Q����\��h�����u�u�%�&�0�>����-���� 9��Z1�\ʴ�1�}�%�6�9�)����I����K��X ��*���g�c�
�g�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����H����@��YN�����&�u�x�u�w�<�(���&����W��h�����%�:�u�u�%�>����	����l��F1��*���
�&�
�y�2�4����K����R��h����u�0�<�_�w�}�W���Y���F��h��*���
�d�d�i�w�u��������\��h_��U���&�2�6�0��	��������F��SN�����%�6�;�!�;�l�G������\��h��D���
�g�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E��Y����T��E�����x�_�u�u�'�.�������� 9��D��*���6�o�%�:�2�.��������V��c1��Gފ�&�
�f�u�/�)��������
U��GךU���0�<�_�u�w�}�W���Y���R��^	�����d�f�i�u��-��������Z��S�����2�6�0�
��.�Eہ�
����F��SN�����;�!�9�d�g�`��������U��W�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�a�}����Ӗ��P��N����u�%�&�2�5�9�E��&����T��E��Oʥ�:�0�&�4��4�(�������@��h��*��u�-�!�:�3����O����l�N�����u�u�u�u�w�}�W�������T9��S1�C���h�}�4�
�8�.�(�������F��h��*���$��
�!�d�;���PӇ����F��*���&�
�#�
�w�}��������U��X�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�f�j�����Ƽ�\��D@��X���u�4�
�<��9�(��N����Z��G��U���'�6�&�}�9�/����I����W9��V
�� ��g�%�y�4��4�(�������@��Q��@���-�!�:�1��(�F��&���F�U�����u�u�u�u�w�}�WϿ�&����Q��_�U��}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ�����]9��D��E���4�
�0�1�1��F݁�K����C9��Y�����e�u�'�;�#�u��������EW��S�����:�1�
� �f�j�(��P����F�R �����0�&�_�_�w�}�ZϿ�&����Q��\����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h-�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�g�w�`�_�������l
��h_��U����
�&�}�w�2����H����F�R �����0�&�_�_�w�}�ZϿ�&����Q��]����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������F��^�����3�
�e�e�'�t�W�������9F�N��U���u�u�u�%�$�:����K���F�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����|�4�1�}�/�)����&����P��G\��U���6�;�!�9�f�m�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6��������� F��D��U���6�&�{�x�]�}�W���
����W��]�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����a�u�h�}�'�>�����ד�[��G1��*���}�u�:�;�8�o�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��X�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�d�;���s���Q��Yd��U���u�u�u�u�w�<�(���&����R��S��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�g�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h\�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�f�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h\�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�a�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h\�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�`�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h]�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�c�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h]�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�l�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h]�U��}�%�6�;�#�1�F��DӇ��p5��D��Bʱ�"�!�u�b�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����I�ƭ�@�������{�x�_�u�w�-��������Q��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��E���h�}�%�6�9�)����H����C9��h��]��1�"�!�u�n�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lR��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����e�1�"�!�w�m�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����������^	�����0�&�u�x�w�}��������W9��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��i�u�4�
��;�������\F��S�����;�!�9�d�f�f�W�������A	��D����u�x�u�%�$�:����M����@��YN�����&�u�x�u�w�<�(���&����U��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��A��i�u�4�
�8�.�(���&���R��d1����u�:�;�:�e�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����l�i�u�4��2����¹��F��h-�����g�u�:�;�8�o�^��Y����]��E����_�u�u�x�w�-��������_��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��Y�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����a�l�i�u�6�����&����F�V��&���8�g�u�:�9�2�E���B����������n�_�u�u�z�}��������lS�������%�:�0�&�w�p�W�������T9��S1�A���&�2�
�'�4�g��������^��1����l�|�u�u�5�:����Y���F�N��U���&�2�7�1�b�i�K������G��Z�����l�d�h�4��2��������F��SN�����8�
�a�'�0�o�N���Y����\��h��*���u�;�u�:��)���&����_��S�����;�!�9�g�g�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������@��1�����0�1�3�
�f��E���	����l��F1��*���
�&�
�y�2�4����J����T��h����u�0�<�_�w�}�W���Y���F��h��*���
�b�u�h��<�(���
����T��N�����<�
�&�$���ف�
������ ��]¼�
�0�0�
��8��������lT��h�Hʴ�
�:�&�
�!��^����Ƣ�GN��G1�����9�d�e�h�2�4����J����T��h�\��u�u�0�1�'�2����s���F������7�1�c�b�6�.��������@H�d��Uʴ�
�<�
�1��j�(�������A	��N�����&�4�
�<��.����&����U��B�����:�1�
� �f�k�(��s���Q��Yd��U���u�u�u�u�w�<�(���&����Q��S��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�w�3�W���Qۃ��G��S[�� ��c�
�g�h�6�����&����O�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����m�4�&�2�w�/����W���F�V�����1�
�m�
�$�4��������C��R������3�8�_�w�}����s���F�N��U���4�
�<�
�3��O���D�έ�l��D��ۊ�u�u�%���.�_�������Q�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����`�4�&�2�w�/����W���F�V�����1�
�l�
�$�4��������C��R������3�8�_�w�}����s���F�N��U���4�
�<�
�3��N���D�έ�l��D��ۊ�u�u�%���.�_������\F��G�U���0�1�%�:�2�.�}�ԜY�����D�����b�g�4�&�0�}����
���l�N��*���
�1�
�e��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��Y���R��X ��*���
�u�u�%������Mӂ��]��Z��N���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�����Y����T��E�����x�_�u�u�'�.��������l��1�����4�&�2�
�%�>�MϮ�������D�����f�l�_�u�w�8��ԜY���F��F��*���
�1�
�c�~�)����Y���F�N�����2�6�0�
��.�F߁�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����l ��hW��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�l�(���&����@��YN�����&�u�x�u�w�<�(���&����l5��D�*���
�e�4�&�0�����CӖ��P�������7�1�c�`�]�}�W������F�N��U´�
�<�
�1��d�^Ϫ���ƹF�N��U���%�&�2�6�2��#���H¹��^9��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���H����^9�������%�:�0�&�w�p�W�������T9��R��!���d�
�&�
�f�<����&����\��E�����%�&�2�7�3�l�A���Y����V��=N��U���u�3�}�%�$�:����H������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���g�3�8�d�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�f�����K����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�f�1�0�F���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:�����3�8�d�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	���&����U��D�����:�u�u�'�4�.�_���
����W��V��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��D��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�a�3�:�l�W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�C�������[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��h�����
�!�`�3�:�l�W�������A	��D�X�ߊu�u�%�&�0�>����-����9��Z1�*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�b�g�u�?�3�}���Y���F�V�����&�$��
�#�h����H�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$����ӓ�@��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�k����H�ƭ�@�������{�x�_�u�w�-��������`2��C_�����d�
�&�<�9�-����Y����V��V�����1�
�b�b�]�}�W������F�N��U´�
�<�
�1��j�@������F�N��U���4�
�<�
�$�,�$����Г�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��X�����`�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����ѓ�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�b�3�8�f���������PF��G�����4�
�<�
�3��F���Y����V��=N��U���u�3�}�%�$�:����H���G��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�c�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*��4�&�2�u�%�>���T���F��h��*���$��
�!�o�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lU��N�����u�u�u�u�w�}��������V��c1��DҊ�&�
�b�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�d�
�$��@��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��Dӊ�&�
�m�4�$�:�W�������K��N�����<�
�&�$����������9��D��*���6�o�%�:�2�.��������W9��Y��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��D��|�!�0�u�w�}�W���Y����C9��P1������&�d�
�$��O��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�Fց�
����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�d�3�:�m�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�\���u�7�2�;�w�}�W�������C9��P1����|�!�0�u�w�}�W���Y����C9��P1������&�d�3�:�m�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�l����I���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���g�
�&�
�n�<����Y����V��C�U���4�
�<�
�$�,�$����֓�@��1�����
�'�6�o�'�2��������T9��S1�B�ߊu�u�0�<�]�}�W���Y���R��^	�����e�|�!�0�w�}�W���Y�����D�����
��&�g��.�(��E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	���&����_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�g��.�(������]F��X�����x�u�u�4��4�(�������@��h��*���4�&�2�
�%�>�MϮ�������D�����a�b�_�u�w�8��ԜY���F��F��*���
�1�
�d�~�)����Y���F�N�����2�6�0�
��.�Eށ�
����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�E݁�
������^	�����0�&�u�x�w�}��������V��c1��G؊�&�
�d�4�$�:�(�������A	��D�����2�7�1�a�`�W�W�������F�N�����4�
�<�
�3��D�������9F�N��U���u�%�&�2�4�8�(���
����U��_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C\�����g�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��\�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�g�
�&��o��������\������}�%�&�2�5�9�C��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���f�3�8�g�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�e�����J����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�g�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�a�1�0�E���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��؊�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�E����ד�@��Y1�����u�'�6�&��-��������W�N�����;�u�u�u�w�4�Wǿ�&����Q��\�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��*���
�u�&�<�9�-����
���9F������6�0�
��$�n����K����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:��ي�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��CZ�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�c�;��������]9��X��U���6�&�}�%�$�:����K���F�U�����u�u�u�<�w�<�(���&����P�����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��h��*���&�<�;�%�8�8����T�����D�����
��&�`�1�0�C���
����C��T�����&�}�%�&�0�?���H���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��C[�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GP��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�c�3�:�h��������\������}�%�&�2�5�9�E��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:��܊�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����l ��hX�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�b�3�8�a�<����&����\��E�����%�&�2�7�3�n�F�ԜY�Ʈ�T��N��U���<�u�4�
�>�����J����[��=N��U���u�u�u�%�$�:����&����GQ��D��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
�ޓ�@�������%�:�0�&�w�p�W�������T9��R��!���m�3�8�b�6�.���������T��]���&�2�7�1�a�e�}���Y����]l�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�%�&�0�>����-����l ��hY��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��CV�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���@����l^��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=�����3�8�m�4�$�:�(�������A	��D�����2�7�1�d�b�t�W�������9F�N��U���}�%�&�2�5�9�F��PӒ��]FǻN��U���u�u�%�&�0�>����-����l ��hV��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��CW�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN���������"�-���N�Փ�lV��1��*��f�%�u�h�]�}�W���Y����u#��u/����� �
�d�
���(���&����D��F�����%�
� �d�f��E��Y���O��[�����u�u�u�'���3���2����F��Y��*���
�
�0�
�c�f�W�������v#��v-�� ���!�g�b�f�2�m�F݁�����9��R�����u�u�u�9���/�������T��R1�����c�f�"�0�w�.����	�Г�F9�� \��G��u�u�d�|�2�.�W���Y�����~ ��-���!�'�
�g���(���&����9F���*������ �'�)�E���J����lW��Q��A���%�u�h�_�w�}�W�������v>��e����a�0�e�'�0�k�Fϩ�����V
��Z�*���d�m�
�g�g�}�W��PӃ��VFǻN��U���'�
������������lU��h^��G���
�a�m�%�l�}�WϿ�����w$��|�����g�b�f�0�g�l�(���H����CU�
NךU���u�u�9����%�������9��1����`�"�0�u�$�1����A����S��h�E���u�d�|�0�$�}�W���Y����A��r+��4��� �%�!�g�`�n����H����lW��1��N���u�4�'����4�������W��1��E���3�
�d�g�'�}�J�ԜY���F��E1��0����:�!� ��l�(���&����T9��N�����&�9�!�%��(�F��&���F�_��U���0�_�u�u�w�}����<����p-��C��*��
�
�
�
�"�l�Oց�J���F��E1��0����:�!� ��l�(܁�&ù��U��_�����h�_�u�u�w�}����<����p-��C��*��
�
�
�
�2��F������@��C��*���d�d�
�g�g�}�W��PӃ��VFǻN��U���'�
������������lU��h^��*���d�e�
�f�]�}�W���&����q'��X�� ���d�
�
�
�����K����Z�=N��U���u�'�
����<���	����Q��h��*���
�c�u�=�9�u��������lW��1��]���h�r�r�u�;�8�}���Y���R��q+��7���:�!� �
�f��(߁�&����T��=N��U���
�����(����K�ѓ�l��hZ�� ��f�
�f�i�w�}�W���YӇ��l ��s,��>���%�!�g�b�2�m�E���������YN�����8�g�3�
�g�j����P���A�R��U���u�u�u�4�%��2���:����C��_��F���e�f�3�
�f�n���Y����A��r+��4��� �%�!�g�`�n����L����W��h�I���u�u�u�u�6�/�1���;����F��C1�B���e�g�'�2�c�o� ���Yە��l��1��*��e�%�}�|�j�z�P������F�N���������8�)����HĹ��V9��1��*��d�%�n�u�w�<����<����x	��G��G���f�0�e�b�1��F���	���l�N��Uʴ�'�����2����&����9��1����l�"�0�u�$�1����&����_��G\��\��r�r�u�9�2�W�W���Y�ƭ�A9��r*��6���!� �
�d���(߁�&����U��=N��U���
�����(����K�ѓ�l��hV�� ��`�
�f�i�w�}�W���YӇ��l ��s,��>���%�!�g�b�d�8�G������� R��_��]���
�8�a�3��l�G���Q���A��N�����u�u�u�u�6�/�1���;����F��C1�B���0�e�b�3��l�@���B�����h(��1���� �%�!�e�j�D���I����V��h�I���u�u�u�u�6�/�1���;����F��C1�B���e�f�'�2�c�m� ���Yە��l��h��D��
�g�e�u�w�l�^ϻ�
��ƹF�N���������"�-���N�֓�lV��R	��C��u�u�4�'���5�������G9�� 1�����d�
� �d�e��D��Y���F���*������ �'�)�E���I����l��hZ�U���;�}�0�
�:�i����J����O�I�\ʰ�&�u�u�u�w�}����?����r%��B����b�f�0�d�n�/���A���F��E1��0����:�!� ��l�(܁�&¹��l ��[�*��i�u�u�u�w�}����7����a4��E��G؊�
�
�0�
�c�}����Q����G��1��*��g�%�}�|�j�z�P������F�N���������2�0�E����ד�V��_�U���4�'������������9��R1��Dي� �d�g�
�d�a�W���Y�����~ ��-���!�'�
�g���(���&����D��F�����%�b�3�
�c�k����P���A�R��U���u�u�u�4�%��2���:����C��_��F���d�d�
� �f�l�(��s���R��q+��7���:�!� �
�f��(���&�ӓ�F9��^��F��u�u�u�u�w�>�(���<����G��h\�*���
�0�
�`�w�5��������CW��Q��@���%�}�|�h�p�z�W������F�N��������:�#�(�(��&����9��h��D��
�f�_�u�w�/�(���=����\��B��D݊�
�
�
�
�"�l�@ׁ�J���9F�N��U���
�����(����K�ѓ�lW��h��*��u�=�;�}�2���������W��G��U��|�0�&�u�w�}�W�������v#��v-�� ���!�g�b�f�2�l����H�ד� ]ǻN���������"�-���N�Փ�lW��h��D��
�f�i�u�w�}�W�������v#��v-�� ���!�g�b�0�f�n����J����[����*���a�'�2�f�e�u�^��^���V
��d��U���u�4�'����4�������W��1��D���3�
�d�m�'�f�W�������v#��v-�� ���!�g�b�f�2�l�D���&����l��S��U���u�u�4�'���5�������G9�� 1�����'�2�a�g� �8�Wǭ�����l��h]�M��u�u�d�|�2�.�W���Y�����h(��1���� �%�!�e�j����K����lU��d��Uʴ�'�����2����&���� 9��1�����d�l�%�u�j�W�W���Y�ƭ�A9��r*��6���!� �
�d���(݁�����F��R �����!�%�
�0��m�C��Y���O��[�����u�u�u�'���3���2����F��Y��*���
�
� �d�n��D�ԜY�ƭ�A9��r*��6���!� �
�d���(ށ�&����V��G]��H�ߊu�u�u�u�%��2���8����G��h\�*���
�
�0�
�`�}����Q����G��h��*��d�e�u�u�f�t����Y���F���*������ �'�)�E���J����lR��B1�Lӊ�f�_�u�u�%��2���8����G��h\�*ي�
�
�
� �f�l�(��E��ƹF�N���������"�-���N�֓�lW��R	��M���=�;�}�0��0�E�������N��S��D���0�&�u�u�w�}�WϿ�����w$��|�����g�b�f�0�f�k����J����F�V��3�����:�!�"��F؁�&����9��h_�E���u�h�_�u�w�}�W���&����q'��X�� ���d�
�
�
������A�ƻ�V�D�����
�0�
�e�f�m�W���H����_��=N��U���u�'�
����<���	����Q��h��*݊� �d�d�
�d�W�W�������v"��t%�����
�d�
�
�����N¹��Z�=N��U���u�'�
����<���	����Q��h_��*���
�c�u�=�9�u��������T9��V��\��r�r�u�9�2�W�W���Y�ƭ�A9��r*��6���!� �
�d���(ށ�����]ǻN���������"�-���N����lV��h��D��
�f�i�u�w�}�W�������]��[�*���=�;�}�0��0�F���&����l��G��U��|�0�&�u�w�}�W�������v#��v-�� ���!�g�b�0�g�m�E�������l�N��������:�#�(�(��&����9��Q��F���%�u�h�_�w�}�W�������v"��t%�����
�d�
�
���(���&����D��F�����%�
� �d�e��E��Y���O��[�����u�u�u�0��0�F߁�����9��d��Uʴ�'�����2����&����V9��1�����f�g�%�u�j�W�W���Y�ƭ�A9��r*��6���!� �
�d���(݁�&����^��@��U¦�9�!�%�
�"�l�E݁�K���F�G�����_�u�u�u�w�8�(���L����U��h����u�'�
����<���	����Q��h^��*ي� �d�g�
�d�a�W���Y�����h(��1���� �%�!�e�j����J�ԓ�V�� ^�����}�0�
�8�f�;�(��K����O�I�\ʰ�&�u�u�u�w�}��������U��_����u�u�4�'���5�������G9�� 1��D���f�3�
�a�o�-�W��s���F�V�����
�#�g�e� �8�Wǭ�����9��h_�G���}�|�h�r�p�}����s���F�V��3�����:�!�"��F؁�&¹��9��P1�E�ߊu�u�'�
���6�������lT��h��*ۊ�
� �d�a��n�K���Y���F��E��0����� �%�#�o�@���H�ד�l��h[�U���;�}�0�
�:�l����J�ԓ�N��S��D���0�&�u�u�w�}�Wϭ�����S��B1�F؊�f�_�u�u�%��2���8����G��h\�*���
�
�
� �f�o�(��E��ƹF�N���������"�-���N����lT��h��*��u�=�;�}�2���������T��F�U���d�|�0�&�w�}�W���Yӕ��l��Z�� ��d�
�f�_�w�}����<����p-��C��*��
�
�
�
��(�F��&���FǻN��U���'�
������������l��h]��*���
�f�u�=�9�u�����ד�F9��\��G��u�u�d�|�2�.�W���Y�����h��D؊� �d�l�
�d�W�W�������l ��h"����
�
�e�3��i�C���Y���F�N����� ���0�:�l�N���H����lQ�������0�
�8�d��8�(��O���F�G�����_�u�u�u�w�/�(���?����\	��\��*ӊ� �g�g�
�d�W�W�������l ��h"����
�
�
� �e�j�(��E��ƹF�N�������!�'��e��������T��N�����&�9�!�%�o�/���N����[�I�����u�u�u�u�w�<��������A��1�����b�b�_�u�w�/�(���?����\	��\��*ي� �g�m�
�d�a�W���Y�����u;��9���'�
�m�0�e�;�(��K����D��F�����%�c�'�2�d�i�_���D����F��D��U���u�u�4�'�9�9�(�������9��P1�L�ߊu�u�'�
�#���������lU��h��G��
�f�i�u�w�}�W�������\��C��*���e�'�2�b�n�*����
����^��h��*��c�e�u�u�f�t����Y���F���*����'��:��o�D�������S��UךU���'�
�!��%�����K�Փ�l ��]�*��i�u�u�u�w�}����,����G��h\�����3�
�f�g�'�}����Q����G�� 1����c�}�|�h�p�z�W������F�N��*�����0�8�f�d��������W��N�����9�
�:�
�8�-�E݁�&Ź��lT��1��U��_�u�u�u�w�1�5���5����^9��1��E���2�b�d�"�2�}��������l��h]�F��u�u�d�|�2�.�W���Y�����h��3����:�
�g�d�h����J�ߓ� ]ǻN�����!��'��8��E���N����R��h�I���u�u�u�u�4��"���<����lW��h��*���
�a�u�=�9�u��������A��_�]���h�r�r�u�;�8�}���Y���R��[�����:�%�g�
�����IŹ��l�N�����
�:�
�:�'�o�(܁�&����T��G]��H�ߊu�u�u�u�;��9�������Q��R1�����b�f�"�0�w�.����	�ѓ�V��X�E���u�d�|�0�$�}�W���Y����_9��y*�����
�m�0�g�1��D���	��ƹF��E�����'��:�
�e�n�N���&����l��S��U���u�u�6�
���2�������l��h��*���u�=�;�}�2����&���� W��^��H��r�u�9�0�]�}�W���Y����_��X�����g�
�
�
�"�o�E߁�J���F��E1��*���
�:�%�g���(߁�I����_��h�I���u�u�u�u�4��"���<����lW��h��*���
�e�u�=�9�u��������A��_�]���h�r�r�u�;�8�}���Y���R��[�����:�%�g�
���(ց�����
9��d��Uʴ�'�9�
�:��2���&����9��Q��L���%�u�h�_�w�}�W�������U��_��]���
�8�d�
�2��F��I���W����ߊu�u�u�u�;��9�������P��R1�����b�`�_�u�w�/�(���?����\	��V��*���
�
� �d�g��D��Y���F���*��f�"�0�u�$�1����O����lU��F�U���d�|�0�&�w�}�W���YӅ��q3��{+�����c�
�
�
�2��@��Y����A��C1�����:�
�m�f�2�m�C���&����l��S��U���u�u�6�
���2�������l��h��*��u�=�;�}�2����&���� W��^��H��r�u�9�0�]�}�W���Y����_��X�����g�
�
�
�����IĹ��l�N�����
�:�
�:�'�o�(܁�&ù��U��\�����h�_�u�u�w�}����I����[����*���d�
�0�
�f�o�G���Y�����RNךU���u�u�9�������&����V9��E��B��_�u�u�'��)�1���5����^��h��*܊� �d�g�
�d�a�W���Y�����u;��9���'�
�c�
������A�ƻ�V�D�����c�'�2�f�c�u�^��^���V
��d��U���u�4�'�9��2�(���	���� 9��1�����l�d�%�n�w�}��������A9��X��M���0�e�b�3��d�B���Y���F�N����� ���0�:�l�N���M����lQ�������0�
�8�d��8�(��O���F�G�����_�u�u�u�w�/�(���?����\	��V��*���
�
� �d�e��D�ԜY�ƭ�A9��h(��*���%�g�
�
���(���H����CU�
NךU���u�u�9�������&����V9��E��M��"�0�u�&�;�)��������P��G��U��|�0�&�u�w�}�W�������T��=N��U���
�!��'��2�(���J����l_��B1�Aӊ�f�i�u�u�w�}�WϽ�&����#��E��Cӊ�
�
�0�
�g�}����Q����G��1����a�}�|�h�p�z�W������F�N�����
�:�
�:�'�o�(܁�&ù��U��Z����u�u�4�'�;���������9��R1��Dڊ� �g�d�
�d�a�W���Y�����u;��9���'�
�c�
������M�ƻ�V�D�����m�'�2�f�`�u�^��^���V
��d��U���u�4�'�9��2�(���	���� 9��1�����e�g�%�n�w�}��������A9��X��M���0�d�d�3��d�D���Y���F�N�����d�d�u�=�9�u��������A��_�]���h�r�r�u�;�8�}���Y���P
��b ��0���8�d�l�0�f�/���J���F��E1��*���
�:�%�g���(ށ�&����
Q��G]��H�ߊu�u�u�u�2��G��������h��D܊�0�
�d�f�g�}�W��PӃ��VFǻN��U���9����#�/�(��&����A��\����u�'�
�!��/�;���&�ޓ�l��hZ�� ��b�
�f�i�w�}�W���YӅ��q3��{+�����c�
�
�
�2��E������@��C��M���2�f�b�}�~�`�P���Y����l�N��Uʴ�'�9�
�:��2���&����9��Q��L���%�n�u�u�6�/��������\��1�����`�3�
�l�c�-�W��s���F�E��D��u�=�;�}�2����&���� W��^��H��r�u�9�0�]�}�W���Y����f(��r����l�0�`�'�0�e�@�ԜY�ƭ�A9��h(��*���%�g�
�
���(���H����CU�
NךU���u�u�9�������&����V9��E��M��"�0�u�&�;�)��������R��G��U��|�0�&�u�w�}�W�������G9��E1�����m�f�0�d�b�;�(��M����9F���*����'��:��e�D���H�ѓ�F9��V��F��u�u�u�u�w�>�(���=����A��W��*ߊ�0�
�f�u�?�3�_���&����9��P1�B���|�h�r�r�w�1��ԜY���F��E1��*���
�:�%�g���(ށ�&����
_��G]�U���4�'�9�
�8�����K˹��V9��1��*��`�%�u�h�]�}�W���Y����f(��r����l�0�b�'�0�e�Nϩ�����V
��Z�*���
�d�g�e�w�}�F�������9F�N��U���
�e�b�_�w�}��������l*��G1�*ي�
�
�
� �e�l�(��E��ƹF�N�������!�'��k�(���&����R��@��U¦�9�!�%�c�%�:�D��Q���A��N�����u�u�u�u�6�/��������\��1�����m�3�
�e�b�-�L���YӇ��l
��q��9���
�c�f�0�g�l�(���K����CU�
NךU���u�u�'�
�#���������l��h]��*���
�l�u�=�9�u��������A��_�]���h�r�r�u�;�8�}���Y���R��[�����:�%�f�
���(ց�����9��d��Uʴ�'�9�
�:��2���&����9��h��G��
�f�i�u�w�}�W�������G9��E1�����c�f�0�e�e�/���Jӑ��]F��R����
� �g�b��o�G���Y�����RNךU���u�u�'�
�#���������l��h]��*���
�l�n�u�w�<����&����	��h]��F���e�d�
� �e�d�(��E��ƹF�N�����!��'��8��A���I�ԓ�l��hV�U���;�}�0�
�:�n�(���K����CT�N��R��u�9�0�_�w�}�W�������l ��h"����
�
�
�
�e�;�(��L����9F���*����'��:��k�D���I����U��_�����h�_�u�u�w�}��������l*��G1�*ي�
�
�0�
�a�}����Q����G�� 1��*��b�%�}�|�j�z�P������F�N�����9�
�:�
�8�-�Dف�&����U��B1�Lӊ�f�_�u�u�%���������C9��h]��*ڊ�
� �g�a��n�K���Y���F��d1��9����!�d�c�c�;�(��O����D��F�����%�m�'�2�d�j�_���D����F��D��U���u�u�4�'�;���������9��R1�����m�d�_�u�w�/�(���?����\	��X��*���
�
� �g�c��D��Y���F���&�����!�d�a�i����J�Г� F��R �����!�%�c�'�0�n�C���P���A�R��U���u�u�u�4�%�1�(���&����lU��1��E���'�2�m�f�]�}�W���&����\��X��F܊�
�
�
�
�"�o�Bځ�J���9F�N��U���
�!��'��2�(���J����lT��R	��B���=�;�}�0��0�Fׁ�����P�N��R��u�9�0�_�w�}�W�������l ��h"����
�
�
�
��(�E��&����F�V�����:�
�:�%�d��(���&ƹ��lT��1��U��_�u�u�u�w��$���:����lW��hZ�� ��a�
�f�"�2�}��������l��h]�G��u�u�d�|�2�.�W���Y�����h��3����:�
�c�2�m�E�������S��N�����9�
�:�
�8�-�Dف�&����9��h\�L���u�h�_�u�w�}�W���&����\��X��F܊�
�
�
�
�2��O������@��C��C���2�f�a�}�~�`�P���Y����l�N��Uʴ�'�9�
�:��2���&����9��Q��A���%�n�u�u�6�/��������\��1�����b�3�
�a�a�-�W��s���F�V�����:�
�:�%�d��(߁�&����T9��N�����&�9�!�%�o�/���N����[�I�����u�u�u�u�w�<����&����	��h]��F���e�c�3�
�c�d���Y����A��C1�����:�
�c�f�2�m�O���&����l��S��U���u�u�4�'�;���������9��1�����2�m�b�"�2�}��������l��h]�G��u�u�d�|�2�.�W���Y��� ��d+��6���!�d�c�a�1��D���	��ƹF��E�����'��:�
�a�n����@����R��h�I���u�u�u�u�6�/��������\��1��E���&�'�2�m�`�*����
����^��h��*��f�e�u�u�f�t����Y���F���*����'��:��k�D���I�ޓ�F9��]��F�ߊu�u�'�
�#���������lU��h_��D���
�`�c�%�w�`�}���Y���R��[�����:�%�f�
���(�������F��R �����!�%�m�'�0�n�@���P���A�R��U���u�u�u�4�%�1�(���&����lU��1��D���3�
�`�l�'�f�W�������G9��E1�����c�f�0�d�f����Mƹ��Z�=N��U���u�'�
�!��/�;���&�Г�l��h\�����g�u�=�;��8�(���Jƹ��lT��1��]���h�r�r�u�;�8�}���Y���R��[�����:�%�f�
���(�������]ǻN�����!��'��8��A����ד� 9��h\�F���u�h�_�u�w�}�W���&����\��X��F܊�
�
�
�
�2��D������@��C��C���
�`�f�%��t�J���^�Ʃ�@�N��U���4�'�9�
�8�����JŹ��V9��\�� ��a�
�f�_�w�}��������l*��G1�*ي�
�
�a�3��k�F���Y���F�N�����9�
�:�
�8�-�Dف�&����A��^����u�&�9�!�'�j����O�ѓ�N��S��D���0�&�u�u�w�}�WϿ�����u	��{��*���f�0�d�d��(�E��&����F�V�����:�
�:�%�d��(���&¹��lT��1��U��_�u�u�u�w����� ����S��R	��G��"�0�u�&�;�)��������Q��G��U��|�0�&�u�w�}�W�������G9��E1�����c�f�0�d�%�:�N��s���R��[�����:�%�f�
���(܁�����9��R�����u�u�u��/�����&�ӓ�V��X����u�&�9�!�'�k����J����O�I�\ʰ�&�u�u�u�w�}��������A9��X��C���0�d�g�'�0�d�F�ԜY�ƭ�A9��h(��*���%�f�
�
���(���K����CU�
NךU���u�u�'�
�#���������lU��h_��*���
�g�u�=�9�u��������A��_�]���h�r�r�u�;�8�}���Y���R��[�����:�%�f�
���(܁�����9��d��Uʴ�'�9�
�:��2���&����9��Q��@���%�u�h�_�w�}�W���*����q��C1�*���
�g�c�"�2�}��������l��h]�G��u�u�d�|�2�.�W���Y�����h��3����:�
�c�2�l�E������� U��N�����9�
�:�
�8�-�Dف�&����9��h\�L���u�h�_�u�w�}�W���&����\��X��F܊�
�
�
�
�2��D������@��C��C���2�f�a�}�~�`�P���Y����l�N��Uʴ�'�9�
�:��2���&����9��Q��@���%�n�u�u�6�/��������\��1�����b�3�
�`�a�-�W��s���F�V�����:�
�:�%�d��(ށ�&����T9��N�����&�9�!�%�o�/���N����[�I�����u�u�u�u�w�<����&����	��h]��F���d�c�3�
�b�d���Y����A��C1�����:�
�c�f�2�l�O���&����l��S��U���u�u�4�'�;���������9��1�����2�l�`�"�2�}��������l��h]�G��u�u�d�|�2�.�W���Y��� ��O=�����
�`�'�2�d�k�L���YӇ��l
��q��9���
�c�f�0�f�d����L�ߓ� F�d��U���u�4�'�9��2�(���	����V9��1�����l�`�"�0�w�.����	�Г�V��Z�E���u�d�|�0�$�}�W���Y����A��C1�����:�
�c�f�2�l�O���&����l��=N��U���
�:�0�!�%��F݁�&����S��G]��H�ߊu�u�u�u�%��2���8����G��hV��D���4�
�0�
�g�n� ���Yے��l_��Q��G���%�}�|�h�p�z�W������F�N��������:�#�(�(���I����W9��P1�L��u�u�4�'�9�9�(�������lU��h��D��
�f�i�u�w�}�W�������\��C��*��
�
�
�0��d�W����ί�]��B1�@܊�g�e�u�u�f�t����Y���F���*���0�!�'�
�f��(���H����CU��N�����;�1�
�0�:�o�E���K����T��h�I���u�u�u�u�6�/����&����lT��h\�� ��`�
�f�"�2�}����&����S��G\��\��r�r�u�9�2�W�W���Y�ƭ�A9��S�����g�g�g�&�%�:�B��s���R��Y��*���8�g�`�<�f�;�(��I����[��C
�����
�0�!�'�"�.����Q����]	��h����`�<�'�2�b�d�W�������V��G1�����9�g�d�|�]�}�W���&����l��Z1�*���1�%�<�3��j�N���Y���F�N�����;�1�
�0�:�e�(ށ�����F��R �����d�a�3�
�`�h����P���A�R��U���u�u�u�4�%�3��������9��E��B��_�u�u�9���;�������l��h��G��
�f�i�u�w�}�W�������l ��h"����
�
�
�0��o�Aϩ�����V
��Z�*���0�
�f�c�g�}�W��PӃ��VFǻN��U���0�
�8�`�����OŹ��l�N��*����'��:��h��������W��N�U���u�u�u�<��<����&����D��F�����%�m�3�
�b�m����P���A�R��U���u�u�u�&�;�)��������R��UךU���9�9�
�:��2���&����U��Y�����h�_�u�u�w�}��������l�������0�
�8�d��(�F��&���F�_��U���0�_�u�u�w�}��������U��X����u�u�6�
�#���������l��h��D��
�f�i�u�w�}�W�������]�� 1��Eʢ�0�u�&�9�#�-�O���&����l��G��U��|�0�&�u�w�}�W���
����^��h��D��
�f�_�u�w�1��������\�� 1��D���
�c�d�%�w�`�}���Y���Z��V ��*݊�
�u�=�;��8�(���H˹��lW��1��]���h�r�r�u�;�8�}���Y���@��C��C���
�c�a�%�l�}�WϽ�&����\��X��Fߊ�
�
� �d�`��F��Y���Z��V �����!�:�
�g�2�k�W������K�d��Uʶ�
�!��'��2�(����֓�F9�� ]��F��u�u�u�u�w�>�(���?����\	��[��*ڊ� �d�b�
�f�*����
����^��h��D��
�g�e�u�w�l�^ϻ�
��ƹF�N�����8�f�
� �f�k�(��s���P
��C1�����:�
�`�0�f�;�(��J����[�N��U���<�
�4� �;�2����&�ԓ�lQ��_��]���
�8�d�
�"�l�G߁�K���F�G�����_�u�u�u�w�8�(���Jǹ��lW��1��N���u�6�;�
�"�l�Bف�K���W�@��U´�'�;�1�
�2�0�E�������lS��S�����;�!�9�g�g�}����[����F�R�����d�3�
�`�d�-�W��[����[�������l�m�h�4��2����������RN��W�ߊu�u�-�!�8�9�(���H����CT�
N��Wʢ�0�u�<�
�>���������A��[�Hʴ�
�:�&�
�!��^ϻ�
���]ǻN�����:�1�
� �f�j�(��E���F��R ��ۊ�0�
�d�u�w�-��������lR�R��U��n�u�u�0�>�>�������� R��N�U��u�=�;�}�%���������W��^1�����l�h�4�
�8�.�(���&����_��^�����u�-�!�:�3����Où��Z�_�����u�<�'�2�c�e�JϿ�&����G9��1�U���0�w�w�_�w�}��������F9��]��G��u�d�u�=�9�u�D�������[��G1�����9�g�g�u�;�8�U���s���U5��r"��!���
�e�
�
�"�o�Cف�J���9F�N��U���
�����(����K�ѓ�l��h_�����f�e�u�=�9�u��������Z9��P1�C���|�h�r�r�w�1��ԜY���F��[1�����<�3�
�f�g�-�L���YӀ��`#��t:����c�3�
�g�o�-�W��s���F�V�����
�#�g�e� �8�WǪ�	����U��W�����|�h�r�r�w�1��ԜY���F��P1�D��u�u�3�
���#���&�Г�F9��X��F��u�u�u�u�w�>�(���?����\	��[��*ۊ�0�
�g�d� �8�Wǽ�&����\��X��Fߊ�
�
�0�
�e�k�G���Y�����RNךU���u�u�'�
�"�d�F���B��� ��b ��;���!�'�
�g�1��@���	�����[�����:�%�g�
������K����F�Q=�����'��:�
�f�;�(��H����[�N��U���<�
��g�2�m� ���Yە��l��V�� ��e�
�g�e�w�}�F�������9F�N��U���
�8�g�
�"�l�Eہ�J���F��h��3����:�
�f�1��A���	���l�N��Uʼ�
��d�0�g�*����
����^��h��D��
�g�e�u�w�l�^ϻ�
��ƹF�N�����8�f�
� �f�i�(��s���U5��R��*��
�
� �g�f��D��Y���F������:�
�:�%�e��(߁�����Q��_��]���
�m�3�
�d�k����P���A�R��U���u�u�u�3���2�������l��h]�C�ߊu�u��!�%�l�F���M����U��h�I���u�u�u�u�4���������C9��h��*���
�g�c�"�2�}����Aù��T9��\��\��r�r�u�9�2�W�W���Y�ƪ�l5��r-�� ���c�'�2�f�e�f�W�������f*��Y!��*���g�3�
�m�f�-�W��s���F�Q=��8���g��!�m��(�F��&����[����*���m�<�3�
�o�h����P���A�R��U���u�u�u�6��)�1���5����S��h_�����g�e�_�u�w�����-����G9��h��D���
�d�i�u��8����Nǹ��lW�� 1��N���u�3�
���o�8���Aǹ��l��h8��*���d�m�
�g�k�}��������E��X�����;�1�%��$�1�(�������
9��N�� ���2�0�}�%�4�3����H˹��u ��UךU����-� ��9�(�(�������g��h��D��
�f�i�u�w�}�W�������l��h�����6�&�
� �f�i�(��������h��G���3�
�b�`�'�u�^��^���V
��d��U���u�&�9�!�'�4����N�ד� ]ǑN��X���'�
� �l�f�>�W�������A	��D�X�ߊu�u�'�
�"�d�F���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�d�y�6�����
����g9��Y�����c�u�9�9��2�(���	����V9��E��F���y�4�
�<��.����&����l ��hW����<�
�&�$����������J��G1�����0�
��&�e�����@�ƭ�l��h�����
�!�
�&��q��������V��c1��Dۊ�&�
�e�u�'�.��������l��1����y�4�
�<��.����&����U��B�����2�6�0�
��.�F݁�
����F��h��*���$��
�!�a�;���UӇ��@��T��*���&�d�
�&��e�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�}�%�6�9�)���������D�����
��&�d��.�(��Y���R��X ��*���<�
�u�u�'�.��������l�� 1����|�:�u�4��2��������F�V�����&�$��
�#�m����@�ƣ�N��h�����:�<�
�u�w�-��������`2��CV�����|�:�u�4��2��������F�V�����&�$��
�#�l����H����AF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�a�u�'��<�(���
����T��N�����<�
�&�$����������O��Y
�����:�&�
�#��}�W�������A9��X��@���e�'�2�f�b�t�W���Q����\��h�����u�u�%�&�0�>����-����l ��hV�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�l�^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����P��D��@���'�}�4�
�8�.�(���&���P
��C1�����:�
�`�0�g�/���L����]�V�����
�:�<�
�w�}��������B9��h��L���8�d�|�u�%�u��������_	��T1�Hʴ�
�<�
�&�&��(���I����lW����U´�
�:�&�
�!��W�������u	��{��*���0�e�'�2�d�h�^���PӒ��]FǻN��U���u�u�'�
�"�d�F���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʲ�%�3�
�l��8�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�:����&����\��S�����;�%�:�0�$�}�Z���YӁ��l ��W�����1�
�&�<�9�-����Y����V��T�����'��:�
�b�8�G�������J��G1�����0�
��&�f�����N�ƭ�l��h�����
�!�
�&��q��������V��c1��Dۊ�&�
�e�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��G1��*��
�%�:�0�k�}��������ET��d��U���u�0�&�3��u��������\��h_��U���&�2�6�0��	���&����V�X�����:�&�
�:�>��W���	����l��F1��*���`�3�8�d�~�2�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��Y�����}�%�6�;�#�1�F��DӅ��_��X�����f�
�
�
�2��E��P����[��=N��U���u�u�u�'��(�N�������VF������!�9�g�e�]�}�W���Y����l�N��U���u�2�%�3��d�(������F��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�2�'�;�(��&����@��YN�����&�u�x�u�w�:����&����CV��D�����:�u�u�'�4�.�_���&����F��h��3����:�
�d�%�:�D��UӀ��K5��N!��*���'�2�f�c�{�<�(���&����l5��D�*���
�b�u�%�$�:����&����G^��D��Yʴ�
�<�
�&�&��(���H����lW�������6�0�
��$�l�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�<�
�&�&��(���A����lW����]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�c�t�W������F�N��Uʲ�%�3�
�l��m�K�������U��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�F�������F��R ��U���u�u�u�u�0�-����@¹��Z�Q=��&����!�`�
�2��E��s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��Uʲ�%�3�
�l��m�K���*����u	��{��*���'�2�f�a�l�}�W���YӃ��VFǻN��U���u�u�'�
�"�d�F���Y���k>��o6��-���������/���!����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���2�%�3�
�n��FϿ�
����C��R��U���u�u�2�%�1��Nށ�H����Z��G��U���'�6�&�}�2��G��Y����u#��u/����� �
�d�
���(�������V����*������ �'�)�E���J����lW��E��F��y�3�
�!��/�;���&�Փ�V��[�U���&�2�6�0��	���&����Q�V�����&�$��
�#�����UӇ��@��T��*���&�d�
�&��m�W���
����@��d:�����3�8�d�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�m�3�8�f�t�W������F�N��Uʲ�%�3�
�l��l�K�������Q��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�B�������F��R ��U���u�u�u�u�0�-����@¹��Z�V��3�����:�!�"��F؁�&����S��R	��G��_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����U��_��D��u�'�
����<���	����Q��h��*���'�2�f�d�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��M���8�b�|�!�2�}�W���Y���F��E�� ��d�%�u�h�1���������C9��h��*��d�_�u�u�w�}����s���F�N�����3�
�l�
�f�a�W͆�!����k>��o6��-���������/��Y���F��Y
�����u�u�0�1�'�2����s���F�	��*���l�`�%�u�$�4�Ϯ�����F�=N��U���
� �l�`�'���������PF��G�����4�
�<�
�$�,�$����ѓ�@��B�����2�6�0�
��.�Fہ�
����F��h��7���!�`�
�0��o�A���*����2��x��Mފ�
�0�
�g�a�W�W�������F�N�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��A�������9F�N��U���u�'�
� �n�h����DӀ��K5��N!��*���'�2�f�c�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Dފ�&�
�f�|�#�8�W���Y���F�	��*���l�`�%�u�j�;�(���5�Ԣ�F��1�����f�b�n�u�w�}�Wϻ�
��ƹF�N��U���'�
� �l�b�-�W��[����k>��o6��-���������/���[���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����3�
�l�
�f�<����Y����V��C�U���2�%�3�
�n��F���
����C��T�����&�}�0�
�g�j�W���
����@��d:�����3�8�d�y�6�����
����g9��Z�����f�u�9�9��2�(���	����V9��E��F��|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��B���8�d�|�u�?�3�}���Y���F�P�����l�
�d�i�w�1��������\��1��E���2�f�d�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�|�!�2�}�W���Y���F��E�� ��`�%�u�h�%�:�F��B���F����ߊu�u�u�u�w�}��������l��S��-���������/���!����k>��o6��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�0�-����@ʹ��P	�������%�:�0�&�w�p�W�������F9��1�����
�&�<�;�'�2�W�������@N��h��*���$��
�!�f�;���UӒ��l^��E��F��y�&�9�!�'�l��������J��R����
�
�0�
�d�i�W���&����
9��E��F��y�&�9�!�'�j��������J��G1�����0�
��&�e�����H���F��P��U���u�u�<�u��<�(���
����T��N�����<�
�&�$����������O��Y
�����:�&�
�#��}�W���&����
9��E��F��|�4�1�}�'�>�����ד�[��R����
�
�0�
�d�k�W���Y������T�����d�e�h�&�;�)��������lU��G��\ʡ�0�u�u�u�w�}�W�������F9��1�����u�h�4�
�8�.�(���&��ƹF�N�����u�}�4�
�8�.�(�������F��h��*���$��
�!�e�;���PӇ��N��h�����#�
�u�u�:��G�������O��Y
�����:�&�
�#��}�W���&����9��E��F��|�4�1�}�'�>�����ד�[��R����
�
�0�
�d�i�W���Yۇ��P	��C1��D��h�&�9�!�'�d��������O��Y
�����:�&�
�#��}�W���&����9��E��F��|�|�!�0�w�}�W���Y�����h��L���:�6�1�u�j�<�(���
����9��=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�Eށ�
����O��_�����u�u�u�u�w�/�(���@�ߓ�C��RN�U���6�;�!�9�b�h�}���Y���V
��d��U���u�u�u�2�'�;�(��&����W�
N��-���w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����
_��N�����u�'�6�&�y�p�}���Y����U��W��E���&�2�
�'�4�g��������_9��h(��*���%�g�
�
��8�(��I�Ư�l
��q��9���
�b�0�d�%�:�D��UӀ��`#��t:�����
�0�
�f�a�}��������B9��h��D���8�g�y�!�'�e�(���&����F��[1�����<�'�2�f�c�q��������l��R	��F��u�0�
�8�e��(���&����F��[1�����<�'�2�f�a�q��������V��c1��G؊�&�
�d�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�e�t����Q����\��h��*���u�0�
�8�e��(���&����F��SN�����;�!�9�d�g�`��������l��R	��F��u�;�u�:��<�(���
����9��
N�����%�e�<�'�0�n�B���P�Ƹ�V�N��U���u�u�2�%�1��Nց�I���U5��r"��!���
�c�'�2�d�o�L���Y�����^��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�e�t����Q����\��h��*���u�8�
�e�%�:�D��PӇ��N��h�����#�
�u�u�2����&����T9��V�����}�%�6�;�#�1�F��Dӕ��l��^��*���
�f�a�u�9�}��������_��N�����!�%�l�<�%�:�D��PӇ��N��h�����#�
�u�u�2����&����T9��X��\ʡ�0�u�u�u�w�}�W�������F9��1��U��6�
�!��%�����L����l��h]�E�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��^��U���;�_�u�u�w�}�W�������l_��h�I���9�9�
�:��2���&����A��\�N���u�u�u�0�$�}�W���Y���F��E�� ��l�%�u�h�u��/���!����k>��o6��-�������u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���T��Q��Lӊ�d�4�&�2�w�/����W���F�P�����l�
�d�4�$�:�(�������A	��D�����
�:�
�:�'�o�(���&���� T��N��*���
�&�$���)�F���������hV�����f�a�y�&�;�)��������lU��B�����8�g�
�
�2��D��Y����G��1�����f�c�y�&�;�)��������lU��B�����2�6�0�
��.�E݁�
����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ԓ�@��G�����4�
�:�&��+�(���Y����V��R	��F��u�;�u�4��2����¹��F��[1�����<�'�2�f�c�t����Q����\��h��*���u�0�
�8�e��(���&����F��SN�����;�!�9�d�g�`��������l��R	��F��u�;�u�4��2����¹��F��[1�����<�'�2�f�a�t�^Ϫ���ƹF�N��U���'�
� �l�n�-�W������]��[�*��u�u�u�u�2�.����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\ʺ�u�}�%�6�9�)���������D�����
��&�g��.�(��Y������T�����d�e�h�&�;�)��������lU��G�����4�
�:�&��+�(���Y����G�� 1�����f�c�|�4�3�3����	����@��A_��U���0�
�8�g������J���O�C��U���u�u�u�u�w�:����&����CW�
N��*����'��:��j��������T��=N��U���u�9�0�_�w�}�W���Y�ƫ�C9��hW�*��i�u�����/���!����k>��o6��-�����n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}��������l*��G1�*���d�c�
�g�k�}��������E��X�����;�1�<�
�>���������A��[�U���;�<�;�1�6�����&����O�=N��U���
� �d�c��o�K�������T��A�����;�<�;�1�>�/���A���F��P ��]���6�;�!�9�d�l�^�ԜY�ƥ�9��h_�A���u�h�&�1�;�:��������F��P ��]���'�2�c�e�w�}��������C9��Y�����d�|�_�u�w��(���K����CT�
N�����2�6�#�6�8�u��������9��P1�M���u�;�<�;�3�<�(���
���� 9��UךU���
�
� �g�n��E��Y����_	��T1�����}�;�<�;�3�4�(���&����M��Y�����4�
�:�&��+�(���B�����E�����'�4�
�0�3�;�(��&���F�
P��*���0�
�y�:�?�/�J���^��ƹF��X��*���3�
�b�f�'�}�Jϸ�&����}"��C��*���3�
�b�e�'�u�D��Hӂ��]��G�U���9�6��d��(�E��&���F��a��*���3�
�e�g�'�u�GϺ�����U�=N��U���
�
�a�3��m�B���Y����l0��1�*���g�f�
�d�e�}�W�������V�=N��U���
�
�`�3��m�G���Y����l0��1�*���g�c�
�d�d�}��������l�N�����d�
� �g�o��F��Y����_T��1��*��b�%�}�f�z�l��������l�N�����d�
� �g�g��C��Y����_T�� 1��*��g�%�}�e�3�*����J��ƹF��X��*���3�
�d�`�'�}�JϮ�/����Q��B1�E؊�d�g�u�u�w�2����I��ƹF��X��*���d�e�
�a�k�}�$���;����v��Z1�*���d�e�
�d�d�}��������l�N�����`�3�
�d�`�-�W��[����[����*���b�3�
�d�b�-�W���	����@��AV��3���9�0�w�w�]�}�W�������U��[�����h�w�w�"�2�}����/����U��Y�����u�%�6�;�#�1�O���PӃ��VF�UךU���:�9�&�
�"�o�Oځ�K���V�@��U¹�6��d�
�"�o�Dځ�M����C9��Y������|�0�&�w�l�L���Yӈ��_��Q��M���%�u�h�w�u�*��������l ��Y�*��h�4�
�:�$��ׁ�?�Ʃ�@�L�U���;�!�=�`�1��F���	���D�������:�
�
�m�1��F���	���R��X ��*���f�e�u�9�2��U�ԜY�Ƣ�G��1��*��d�%�u�h�u�� ���Yۊ��l0��1��*��e�%�u�u�'�>��������O��[��W���_�u�u�:�%�.�(���K����CT�
N��Wʢ�0�u�9�6��l�(���K����CW������!�9�g�
�~�8����I��ƹF��h^�D���<�3�
�m�f�-�W��s���F�V�����
�#�f�e� �8�WǪ�	����U��^�����|�h�r�r�w�1��ԜY���F��T1��D؊� �d�d�
�f�W�W���&����_��1��*��b�%�u�h���"���7����V��\�� ��e�
�d�f�w�2����J�����hV�����
�m�l�%�~�W�W���&����_��h��D��
�f�i�u�6�����&����lV���*��� �d�e�
�c�f�W���	����9��h��G��
�d�i�u���;���6����9��P1�G��u�u�%��;��A���&����l��S�����
�:�
�:�'�o�(���&���� T��d��Uʥ��9�
�b�1��F���	�����[�����:�%�g�
������K����F�G�����
� �g�g��n�K���Y���F��E��0����� �%�#�o�@����֓�9��P1�E���=�;�}�8��m����J����O�I�\ʰ�&�u�u�u�w�}����<����|��^�����g�m�%�n�w�}����K����l��V�����
� �d�a��n�K���Y���F��G1�����9�d�
�e�w�5��������Z9��_�� ��g�
�g�e�w�}�F�������9F�N��U���6�;�!�9�f��G��Y����V��h��*���d�g�
�f�k�}�W���Y����C9��Y����
�e�e�"�2�}��������lU��Q��B���%�}�|�h�p�z�W������F�N��*���&�
�#�`�c�m�L���Yӕ��l��^�� ��c�
�f�i�w�}�W���YӇ��P	��C1��F؊�u�=�;�}�2���������^��F�U���d�|�0�&�w�}�W���YӇ��l ��s,��>���%�!�g�b�2�m�F�������
V��N�����!�%�d�3��n�C���Y���F�N���������8�)����HĹ��9��1�����e�"�0�u�$�1����&����_��G\��\��r�r�u�9�2�W�W���Y�ƭ�l��D�����e�_�u�u�2����&����lT��1��U��}�8�
� �e�n�(���Ƹ�C9��1�����4�
�
� �e�k�(��B�����h��Dۊ�
�:�
� �e�k�(��E����V
��Z�*��� �g�f�
�e�%�Ͽ�&����G9��1�N���u�&�9�!�'�o����J�ԓ� F�d��U���u�4�'����4�������W��R1��F���'�2�`�e� �8�Wǭ�����9��h_�M���}�|�h�r�p�}����s���F�D�����d�3�
�f�c�-�L���Yӕ��l��\��*���g�g�
�f�k�}�W���Y����A��r+��4��� �%�!�g�`�n����Hƹ��T9��^�����}�0�
�8�f��(���&����V�
N��R���9�0�_�u�w�}�W�������l ��]�*��_�u�u�0��0�F܁�����9��R�����u�u�u�%�4�3����J����D��F�����%�
� �d�n��E��Y���O��[�����u�u�u�'���3���2����F��Y��*ۊ�
�
�0�
�c�f�W���
����^��h��D��
�f�i�u�w�}�W�������v#��v-�� ���!�g�b�0�f�o�E���������YN�����8�m�3�
�d�e����P���A�R��U���u�u�u�&�;�)��������^��UךU���0�
�8�d��(�F��&���FǻN��U���%�6�;�!�;�n�(������@��C��*���d�e�
�g�g�}�W��PӃ��VFǻN��U���'�
������������l��h_��*���
�`�n�u�w�.����	�Г�F9�� \��G��u�d�u�=�9�u����N����R��h�Hʴ�
�:�&�
�!��^ϻ�
���]ǻN�����8�d�
� �f�e�(��E���F��R �����l�
� �d�a��F������]��[��G���9�0�w�w�]�}�W���&����9��h_�E���u�h�w�w� �8�WǪ�	����U��X�����u�%�6�;�#�1�E��Y����D��d��Uʦ�9�!�%�m�>�9��������lT��1��U��}�8�
�l�1��F���	�ƣ���h��Dۊ�
� �g�f��o�L���Yӕ��l��V��*���g�`�
�g�k�}��������l��R�����3�
�g�`�'�}����	����@��A_��\�ߊu�u�0�
�:�l�(���H����CU�
NךU���u�u�;��>�.�C���Kӑ��]F��R����
� �d�b��o�G���Y�����RNךU���u�u�;��>�.�C���O���F��[1�����<�3�
�g�`�-�W��Q����U��B1�Eӊ�g�-�'�4��2����¹��l�N�����%�
� �d�e��E��Y���D��F����
� �d�l��l�JϿ�&����G9��1�U���0�w�w�_�w�}�����ד�l ��Y�*��i�u�!�%�>�4����&����l��O�����:�&�
�#��t�}���Y����G��1��*���a�%�u�h�]�}�W���Y����R��hZ��*���=�;�}�0��0�F؁�����9��^��H��r�u�9�0�]�}�W���Y����G��1��*���m�%�n�u�w�.����	�֓�l ��\�*��i�u�&�9�#�-�O�������W��N��ʦ�9�!�%�l�>�;�(��N����l�N�����%�d�3�
�b�e����D���F�N��*���;�
�
�
�w�5��������CW��Q��A���%�}�|�h�p�z�W������F�N��*���;�
�
�
�l�}�Wϭ�����W��h��G��
�f�i�u�w�}�W�������v#��v-�� ���!�g�b�f�2�m�Fځ�����V��_��]���
�8�g�
��8�(��M���F�G�����_�u�u�u�w�8�(���H����U��\����u�u�&�9�#�-�E���&����l��S��U���u�u�<�
�6�3�(ہ�&�ƻ�V�D�����b�3�
�a�a�-�_���D����F��D��U���u�u�&�9�#�-�F���&����l��=N��U���
�8�g�
�"�l�@ׁ�J���9F�N��U����;�0�b�2�o� ���Yە��l��X�� ��b�
�g�e�w�}�F�������9F�N��U����;�0�b�2�k�}���Y����G��1��*���a�%�u�h�]�}�W���Y����R��hY��*���=�;�}�0��0�F؁�����9��^��H��r�u�9�0�]�}�W���Y����G��1��*���m�%�n�u�w�.����	�ӓ�F9��V��F��u�u�u�u�w�4�(�������V9��@��U¦�9�!�%�c�1��C���	����[�I�����u�u�u�u�w�4�(�������V9��=N��U���
�8�g�
�"�l�Gہ�J���9F�N��U����;�0�b�2�h� ���Yە��l��Y�� ��m�
�g�e�w�}�F�������9F�N��U���
�8�g�
�"�l�Nׁ�J���F��[1�����3�
�c�m�'�}�J�ԜY���F��h>��G���d�"�0�u�$�1����O����R��h�E���u�d�|�0�$�}�W���Y����]9��h\��*��u�u�&�9�#�-�O���&����l��S��U���u�u�<�
��o���������h��D݊� �d�m�
�e�m�W���H����_��=N��U���u�0�
�8�e����H˹��l�N�����%�m�<�3��o�B���Y���G��W�� ��b�
�g�4�3�.����	�ד�l��h��G��
�g�n�u�w�.����	�ߓ�F9��V��F��u�u�u�u�w�4�(���H������YN�����8�d�
� �f�j�(��I���W����ߊu�u�u�u�%���������W��1�����a�`�_�u�w�8�(���Kʹ��U��V�����h�}�8�
�a�;�(��H����R��D�����m�<�3�
�e�h����s���@��C��*���d�l�
�g�k�}�F������G��Z�����l�d�h�4��2����������RN��W�ߊu�u�0�
�:�o����&����l��S�����d�d�<�<�>�;�(��N����R��D�����
�
� �d�b��E��Y����V
��Z�*���d�a�
�f�k�}�W���Y����A��X
�����
�d�
�
��8�(��Y����N��[1�����3�
�a�c�'�u�^��^���V
��d��U���u�&�9�!�'�d����O�ޓ� ]ǻN�����8�f�
�
�"�o�C߁�J���9F�N��U���
�����(����K�ѓ�l��h_�����f�e�u�=�9�u��������Z9��P1�C���|�h�r�r�w�1��ԜY���F��[1�����<�3�
�f�c�-�L���Yӕ��l��_�� ��c�
�d�i�w�m�I���4����_%��C��*���0�a�u�!�2�.�I��P���F��[1�����3�
�c�e�'�}�J���D͏��~��V�����9�d�
�
�{�2����D���]ǻN�����8�f�
� �f�k�(��E��ƹF�N�����8�f�
� �f�k�(��������h��D܊� �d�b�
�e�m�W���H����_��=N��U���u�0�
�8�d����Où��l�N�����%�g�3�
�a�k����D������z�����;�'�9�d���[ϱ�����A�UךU���0�
�8�f��(�F��&���FǻN��U���0�
�8�f��(�F��&����[����*���d�
� �d�o��E��Y���O��[�����u�u�u�0��0�Dށ�����9��d��Uʦ�9�!�%�f�1��A���	���l�N��Uʼ�
�4� �9�8�)����K������YN�����8�d�
� �f�j�(��I���W����ߊu�u�u�u�9�����:����\
��1��F�ߊu�u�0�
�:�n�(���H����CU�
NךU���u�u�;��9�<�4�������9��N�����&�9�!�%�`�;�(��O����O�I�\ʰ�&�u�u�u�w�}��������l ��X�*��_�u�u�0��0�Dځ�����
9��R��W���"�0�u�!�'�l�D���&����l��
N��*���&�
�#�
�~�8����I��ƹF��R����
� �g�l��o�K���H�ƻ�V�C��D���3�
�`�`�'�}�W�������l
��h\�����u�e�n�u�w�.����	�ѓ�F9��Y��G��u�d�u�=�9�u����I����lT��1��U���%�6�;�!�;�o�G������D��N�����!�%�b�<�1��E���	���N��G1�*���g�e�
�g�6�9��������l��B1�@ۊ�g�n�u�u�$�1����&���� U��G]��H�ߊu�u�u�u�'�>��������F��R �����!�%�
� �f�d�(��I���W����ߊu�u�u�u�%��2���8����G��h\�*���
�
�
�0��e�L���Yӕ��l��_��*���g�`�
�f�k�}�W���Y����C9��Y����
��e�e�g�*����
����^��h�����f�m�e�u�w�l�^ϻ�
��ƹF�N��&���'�d�d�g�c�;�(��N����9F���*���a�3�
�d�g�-�W��[����[����*���'�2�g�l�w�}��������ET��N�����e�n�u�u�$�1����I����F9��W��F��u�u�u�u�w�;�(���¹��9��Q��F���%�u�=�;��8�(���Kù��A��]�]���h�r�r�u�;�8�}���Y���@��C��D���3�
�f�g�'�f�W���
����^��h�� ��c�
�f�i�w�}�W���YӅ��_��X�����g�
�
�
�2��E��������h��Gӊ�
�0�
�f�g�m�W���H����_��=N��U���u�0�
�8�b��(���K����CU��N�����!�%�
� �f�i�(��E��ƹF�N���������"�-���N����lT��h��*��u�=�;�}�2���������^��F�U���d�|�0�&�w�}�W���Yӕ��l��1��*��c�%�n�u�w�.����	Ź��lW��1��U��w�w�"�0�w�)���&����_��G_��U���6�;�!�9�e�o�W�������l�N�����%�
�
� �f�k�(��E���F��R �������g��#�e�(�������V9��h_�D���u�u�%�6�9�)���&����F��D��E��u�u�&�9�#�-�(���H����CU�
NךU���u�u�'�
���6�������lT��h��*ي�
�0�
�b�w�5��������CP��B1�Lފ�g�e�u�u�f�t����Y���F������!�9�f�
�l�}�Wϭ�����9��Q��M���%�u�h�w�u�*��������f*��Y!��*���<�
�%�,�2�;�(��H����F��h�����#�`�a�e�w�1����[���F��[1��Ҋ� �d�e�
�e�a�W��Y����N��G1�*���d�l�
�d�j�<�(���
����9�������w�_�u�u�2���������^��h�I���&�9�!�%�����O����	��D�����
�
� �d�a��E��Y����V
��Z�����f�a�%�u�j�W�W���Y�ƭ�A9��r*��6���!� �
�d���(܁�&����Q��@��U¦�9�!�%�
�"�l�Gׁ�K���F�G�����_�u�u�u�w�8�(���N����U��h����u�0�
�8��(�F��&���F�N�����!�%�l�
�2��N��DӇ��P	��C1��G��u�9�0�w�u�W�W�������C9��Q��B���%�u�h�_�w�}�W�������Z9��Q��B���%�u�=�;��0�(���&����lW�� 1��]���h�r�r�u�;�8�}���Y���R��X ��*���`�a�e�_�w�}����I����lT��1��U��<�
�0�
�a�u�W���Y����G	�UךU���8�
�e�
�"�o�Gځ�H���ZU��R	��B���u�u�u�:�9�2�G��Y����^��_��*���d�l�
�g�k�}�F������@��R
��&��� ��;� ��i��������9��h_�B���|�i�&�2�2�u��������EW��G�����u�e�n�u�w�)���@����\��Y1�����e�d�%�u�j�u����&�ԓ�l ��^�*��4�1�!�%�>�4�(�������9��UךU���8�
�g�
�2�2��������V��h�I���!�%�<�<���E���&����l��V �����<�<�
�
�"�o�N߁�K��ƹF��Z��Gي�0�:�2�;�>�;�(��H����[�C�����
�
�f�3��l�N���Y����G��^1��*��� �g�g�
�e�f�W������� W��h��*���d�f�
�g�k�}�F������_	��a1��*��f�%�u�u�'�>�����ޓ�uO��[��W���_�u�u�8��d����A�ӓ�F�F�����3�
�b�f�'�}�Ϫ�	����l��B1�Lӊ�g�n�u�u�#�-�A߁�����
9��R�����u�u�u�%�4�3����A����D��F�����3�
�b�f�'�u�^��^���V
��d��U���u�4�
�:�$��ׁ�B�����hX�����m�d�%�u�j�W�W���Y�Ƹ�C9��h��D��
�f�"�0�w�)���&����V��G\��\��r�r�u�9�2�W�W���Y�Ƹ�C9��h��D��
�d�_�u�w�0�(�������
R��N�U¡�%�<�<�<�d����K����	��Y����� �d�m�
�e�f�W�������9��h\�F���u�h�}�8��o����J����R��P�����l�
�g�n�w�}����Oƹ��lT��1��U��}�:�'�&��(�E��&����AF��C��@���
�d�b�%�~�W�W�������l ��_�*��i�u�;�!�?�k����H�ד�F�� �����
� �g�`��o�L���YӒ��lP��Q��D���%�u�h�}�:��B���&����l��V �����c�
� �g�a��E��Y����^��1��*��l�%�u�h��0�(�������U��N��ʲ�%�3�
�l��o�L���YӒ��lQ��Q��D���%�u�h�}�8�/�؁�����9�������=�b�3�
�f�h����s���G�� _�� ��e�
�g�i�w�)���&����_��G\�����8�
�`�3��l�N���P���F��G1�*���d�e�
�%�8�8�K���	����@��A[��N���u�!�%�b��(�F��&���F��h=��0��� �
�c�'�0�n�E��Y����^��1��*��f�%�u�h�4���������C9��h��*���
�g�c�_�w�}����J����T��h�I���!�%�b�
�"�o�G܁�KӇ����hY�����e�f�%�|�]�}�W���&�ғ�F9��[��G��u�!�%�b��(�E��&����]��Z��C���
�d�b�%�~�W�W�������l ��^�*���:�0�i�u�'�>�����ӓ�l�N����
� �d�e��m�K���*����v%��B��C���2�f�g�n�w�}����Nƹ��lW�� 1��U��6�
�!��%�����N����l��h]�B�ߊu�u�8�
�a�;�(��H����[�C��Bފ� �g�d�
�e�<�Ϫ�	����U��^�����_�u�u�8��e����J�Г�F�F����
�0�
�f�`�<�Ϲ�	����
_��G\����u�8�
�l�1��G�������VF������!�9�`�a�]�}�W���&�ߓ�F9��_��E��u��������&���� U��d��Uʡ�%�b�
� �f�l�(��E�Ư�l
��q��9���
�b�0�d�%�:�D��B�����hV�����g�b�%�u�j�u����H����T��h����!�%�b�
�"�l�Fށ�K��ƹF��Z��C���3�
�m�l�'�}�J�������l ��V�*��s�%�e�g���(���H����CU�=N��U���
�a�3�
�g�o����Dӏ��V��V��U���u�:�;�:�g�f�W�������9��h_�C���u�h�4�'�9�9�(�������l��R	��D���u�u�u�:�9�2�G��Y����^��1��*��e�%�u�h�>�����H����F��S�����|�_�u�u�:��@���&����l��S��9���
�:�
�:�'�.����@���K�
�����e�n�u�u�#�-�Nց�����9��R�������g��#�e�(�������lT��B1�M݊�g�m�x�d�3�*����P���F��G1��*��f�%�u�h��0�(��&����A��h�� ��l�
�g�:�w�0�(��&����A��h�� ��f�
�g�n�w�}��������Q��h�I���d�u�=�;��4��������f*��Y!��*���<�
�-�
�����AĹ��F�D�����%�6�;�!�;�l�(���PӃ��VF�UךU���8�
�
�g�>�;�(��@����[�L�����}�:�
�
�d�;�(��L����F��h�����#�
��u�;�8�U���s���G��^1��*���g�3�
�e�c�-�W��[����[����*���`�3�
�e�g�-�W���	����@��AV��3���9�0�w�w�]�}�W���&����l��B1�@ߊ�g�i�u�e�w�5��������R��B1�Aߊ�d�h�4�
�8�.�(���J���V
��L�N���u�!�%�<�>��(�������_��N�U��u�=�;�}�8��(�������S��N�����:�&�
�#���W�������l�N�����<�
�
� �e�d�(��E���F��R ������d�
� �e�e�(��DӇ��P	��C1��Gي�|�0�&�u�f�f�W�������l��^1��*��`�%�u�h�u�� ���Yۊ��l0��1��*��`�%�u�u�'�>��������O��[��W���_�u�u�8���(���H����Q��h�I���d�u�=�;��2�(���K����Q��h�Hʴ�
�:�&�
�!�n�G������D��N�����<�<�<�3��j�@���Y���D��_��]���
�
� �d�g��C������]��[��E���9�0�w�w�]�3�W������