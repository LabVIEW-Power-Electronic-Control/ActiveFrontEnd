-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�M���� ^��1��@���3�`�d�m��<�W���s���T��E�����u�u�u�u�w�8�(������	F��E��U��w�9�6�w�w�}�W���Y�����S��U���o�<�!�2�%�g�W��Y���F�N��U���1�=�u�u�m�4�������]�N��U���u�u�8�8�$�'�W���Cӏ��V��T��G���u�|�u�u�w�-����s���F�N����u�u�o�<�w�)�(�������P�������d�1�"�!�w�t�W���Y���F��R^��U���u�u�;�&�3�1����Y���F�N��E���u�u�u�u�"�}��������E��X�����=�d�1�"�#�}�^�ԜY���F�V
��D���u�o�<�u�#�����&����\��@����1�"�!�u�~�}�W���Y�����N��U���u�;�&�1�;�:����Y���F�
�U���u�u�u�;�$�9��������G	��S�����u�:�;�:�g�f�}���Y���F��N��U���o�<�u�!��2���s���F�N�����u�u�u�u�9�.�������F�U�����0�!�!�n�]�W��������A��C��ʸ�a�c��m���(ځ�����^��h��U���_�&�2�4�w�9�߁�����@��[�����6�:�}�"�3�5�FϺ�����O��=��ʸ�8�4�'�,�>�}����Y����\F��Z1�����|�:�u�!��2��������N��^
��X���:�;�:�e�l�W����Ӑ��Z��RN����8�8�4�'�.�W����������h�����0�o�&�'�9�f�}�������VF��Y1�����9�u�3�'�:�g��������Z�U�����8�n�4�!�>�(�Ϭ�����_������_�!�'�7�#�}��������\ ��V��U���<�7�0�<�w�8�(������G��B��0������
���#���+����r*������_�7�2�;�]�W���� ����V��P����u�'�6�&�w�<���Y����ZǻN��U���'�
�8�u�j�<���s�˿�]��D�����&�4�0�:�1�}�W�������|(��~ ��2���4�1�e�u�w�8�(������G��=N��U���u�u�4�1�g�)���Yۉ��V��
P��E���_�u�u�u�;�8�}���Y���F��S
��*���u�h�4�1�g�W�W���Y����Z ��C�����&�&�!�4�$�<����s����C��R����8�8�'�
�4�8���Y����V����\���7�2�;�_�w�}��������V��V �����h�r�r�u�?�3�W���Y����UF��R^��U��|�!�0�u�w�}�W���Y����F���]��������<�������FǻN��U���;�u�3�_�w�}�������WF��X���ߠ_�
�0�:�.�<����&����A	��D�����u�_�0�<�w�}�WϷ�Yۅ����Y�����9�u�u�d�~�)��ԜY���F��F��D��r�r�u�=�9�W�W���Y���F��F��D��r�r�u�=�9�W�W���Y���F�N����
����u����P������d��U���u�u�u�0�3�4�L���Y����������u�;�u�3�]�3�W�������9l��Y
����_��7�4�.��2������v#��D�����6�d�c�{�;�f�}�������uR��/����3�`�7�3�b�l�O���
�����R��U�ߊu�u�u�u�6�<����Y�ƅ�g#��eN�U��_�u�u�u�w�9����+����\��y:��0���h�g�_�u�w�}�W�������Z��T��;����u�h�d�l�}�WϮ����F�N�����!�o��u���8���B���F���U���������}���Y���R��R��U���������!���6�΍�W��D9�����u�u����m�L���Y�����T��;ʆ�����]�}�W���Y���)��=��*����
�����������W��x9��:��n�u�u�u�w�<����
����z(��c*��:���
�����9��������F��s!��!���|�_�u�u�w�}����Y����g"��x)��N���u�u�u�"�f�g�>���-����t/��=N��U���u�d�o��w�	�(���0����p2��*�����!�u�u�u���8��P���WF��C��N���'�=�!�6�"�8����Y����uR��/����3�`�7�3�b�l�O���
�����G������e�l�f�1�m��������lW��1��ʼ�_�u�u�u�w�2����Y���F�N�����u������4�ԜY���F�N����o��u����>���<����l�N��U���u�6�e�o��}�#���6����9F�N��U���u�e�o����3���>����v%��eUךU���u�u�u�u�3�/�W���7ӵ��l*��~-��0����_�u�u�w�}�W�������z(��c*��:���n�u�u�u�w�}�WϺ�Y�ƅ�5��h"��<������_�w�}�W���Y�ƻ�F��~ ��!�����|�_�w�}��������V��=dװ���;�u�u�8�c�k�6���&ù��9��Q1��D��
�4�
�u�w�>��������uR��/����3�`�7�3�b�l�Oہ����F��E�����_�u�u�u�w�1�W�������F�N�����e�h�u�1�%�.�G�ԜY���F��N��U���y�u�u�u�w�,�W�����ƹF�N�����u�k�4�1�2�.�[���Y�����S���_�u�u�u�w�l�J���H���F�N��D��u�0�|�_�2�9��������F��=d�