-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�a�c��m���(�����A�=N��U���6�>�o��w�	�(���0��ƹF��G1�����u��
���L���YӇ��@��CN�<����
���l�}�WϿ�&����\��b:��!�����n�u�w�<�(�������f2��c*��:���n�u�u�4��8����Y����`2��{!��6�ߊu�u�;���<����&����	F��=��*����
����u�FϺ�����O��N������'�;�0�n�8�F��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����E����o��u����>��Y����]9��{	�����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���)����Z��1��D���u��
���(���-��� W��X����n�u�u�<��)����&ù��F��~ ��!�����
����_������\F��d��Uʼ�
�'�1�-�2�)��������	F��=��*����
����u�FϺ�����O��N������`�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�������/��d:��9�������w�n�W������]ǻN�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W�������G��h_��U���u��
����2���+������Y��E��u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�V�����;�f�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������z(��c*��:���u�n�0�1�]�W��������A��R��U���8�a�c��o��(���Iӏ��9F������!�4�
�:�$�����&����`2��{!��6��u�d�n�u�w�>�����ƭ�l��D�����
�u�u����>���D����l�N�����;�u�%���)�(���&����`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�E��w�_�u�u�8�.��������l��h��*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V�=N��U���&�4�!�4��	��������\��c*��:���
�����d��������\�^�E��e�e�e�e�g�m�G��Y����\��V ������&�`�3�:�i�Mύ�=����z%��r-��'���l�1�"�!�w�t�M���I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�����`�o�����4���:����W��S�����|�o�u�e�g�m�G��I����V��L�U���6�;�!�;�w�-�$���Ĺ��^9��N��1��������}�F�������V�S��E��e�e�e�e�g�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�e�e�w�]�}�W���
������d:��ӊ�&�
�u�u���8���&����|4�W�����:�e�u�h�u�m�G��I����V��^�W�ߊu�u�:�&�6�)����-����9��Z1�Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�l�G��I����l�N�����;�u�%���)�F�������	F��s1��2������u�f�}�������	[�^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�g�3�:�l�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��e�e�w�_�w�}��������C9��h��F���8�d�u�u���8���&����|4�W�����:�e�u�h�u�m�G��H����V��^�W�ߊu�u�:�&�6�)����-����9��Z1�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����]ǻN�����4�!�4�
��.�Fځ�
����\��c*��:���
�����d��������\�^�E��e�e�e�e�g�m�G��Y����\��V ������&�d�
�$��B��*����|!��h8��!���}�l�1�"�#�}�^��Y����W��^�E��e�e�e�n�w�}��������R��c1��D݊�&�
�c�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��^�E��u�u�6�;�#�3�W���*����^��D��B��������4���Y����W	��C��\��u�e�d�e�g�m�G��I����D��N�����!�;�u�%����������F��d:��9�������w�l�W������F��L�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�e�1�0�F���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�e�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�d�d�o���;���:����g)��^�����:�e�u�h�u��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������rF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EU��tN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��_�E��u�u�6�;�#�3�W�������l
��1��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�D��n�u�u�6�9�)����	����@��A]��D���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�e�e�e�e�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�F��I����V��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�
�#�g�`�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�l�F��Y����\��V �����:�&�
�#�e�l�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(ܘ�I����\��c*��:���
�����l��������\�^�D��d�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EU��+��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�D���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Nӂ��]��G��H���e�e�e�e�l�}�WϽ�����GF��h�����#�f�e�o���;���:����g)��\����!�u�|�o�w�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*��e�o�����4���:����W��S�����|�o�u�d�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���L����F��d:��9�������w�l�W������F��L�E��e�e�e�e�g�f�W�������R��V�����
�#�
��m��3���>����v%��eN��U���;�:�e�u�j��F��H���9F������!�4�
�:�$�����L���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����d�
�e�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��L�U���6�;�!�;�w�-��������9��N�&���������W��Y����G	�N�U��e�d�e�e�g�m�G��Y����\��V �����:�&�
�#�g�m�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����V��UךU���:�&�4�!�6�����&����lU��q(��U���
���
��	�%���Nӂ��]��G��H���d�d�d�d�f�l�F��H��ƹF��X �����4�
�:�&��+�O���Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��d�d�d�w�]�}�W���
������T�����d�
�u�u���8���&����|4�Y�����:�e�u�h�u�m�G��I����V��_�����u�:�&�4�#�<�(���
���� T��q-�E��o������!���6���F��@ ��U���o�u�e�d�f�l�F��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�d�w�]�}�W���
������T�����`�`�o����0���/����aF�
�����e�u�h�w�g�m�U�ԜY�Ư�]��Y�����;�!�9�`�f�g�$���5����l0��c!��]���:�;�:�e�w�`�U��I����F�T�����u�%�6�;�#�1�B��Cӵ��l*��~-��0����}�u�:�9�2�G���D����V��d��Uʶ�;�!�;�u�'�>�����ӓ�\��c*��:���
�����}�������	[�^�E��_�u�u�<�9�1����*����\��c*��:���
�����d��������\�^�E��e�e�e�e�g�m�F��Y����G��U��U���
�;�:�<�0�g������ƹF��C�����u�&�
�;�8�4�ϱ�Y����`9��ZN����4�u�&�w�8�8�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������\��x!��4��u�u�&�2�6�}����<����x	��G��F݊�
�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W���������q+��7���:�!� �
�`�m���Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������2�%�3�
�d��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���
����@��d:��ي�&�
�u�u���8���B�����Y�����<�
�1�
�o�g�5���<����F�D�����%�&�2�6�2��#���N����lP�=��*����n�u�u�$�:����	����l��hY�Oʗ����_�w�}����Ӂ��l ��]�����u��
����2���+������Y��E��u�u�&�2�6�}����N����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���&���� F��d:��9����_�u�u�>�3�Ͽ�&����Q��V��U�����n�u�w�.����Y����Q��N��1��������}�D�������V�=N��U���;�9�4�
�>�����*����V��D��U����
���l�}�Wϭ�����R��^	�����m�o�����}���Y����R
��G1�����0�
��&�f�����L����g"��x)��N���u�&�2�4�w�-��������P�,��9���n�u�u�&�0�<�W�������lR��R�����
� �m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����P
��r+��4��� �%�!�f���(ށ�����l��N��1��������}�D�������V�=N��U���;�9�3�
���E�������9��h]�*��o������!���6���F��@ ��U���_�u�u�<�9�1����4����])��hV��G���2�d�`�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����A��\�U����
�����#���Q�ƨ�D��^����u�<�;�9�1��:���K����lP��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������f*��Y!��*���g�'�2�d�a�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h=��0��� �
�a�
�"�k�G���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�������� ��i�(���&����\��c*��:���
�����l��������l�N�����u�%�&�2�4�8�(���
�ӓ�@��T��!�����n�u�w�.����Y����Z��S
��F���u����l�}�Wϭ�����R��^	������
�!�d�1�0�F���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�)���&����
U��N�&���������W������\F��d��Uʦ�2�4�u�8��j����H����	F��s1��2������u�g�9� ���Y����F�D�����8�
�f�3��m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
�0�
�g�o�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��D���3�
�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��D���'�2�d�e�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*��� �m�d�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���0�
�f�e�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G\�����
�`�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G\�����2�d�d�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��Y��*���m�`�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��Y��*���
�f�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����f(��r����
�
�
� �n�o����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*�����0�8�e��(݁�����^�=��*����
����u�FϺ�����O��N�����4�u�%�&�0�>����-����9��Z1�U����
���l�}�Wϭ�����R��^	�����b�u�u����L���Yӕ��]��Q=��8���,� �
� �#�-���&����U��T��!�����
����_������\F��d��Uʦ�2�4�u�%�$�:����&����GW��Q��D���u��
���f�W���
����_F��h��*���
�m�u�u���6��Y����Z��[N��*����� �
�o�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����%�&�2�6�2��#���Hǹ��^9��T��!�����n�u�w�.����Y����Z��S
��L���u����l�}�Wϭ�����Q	��h�����
�m�3�
�g�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T���������!�a��8�(��L����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$����������F��d:��9����_�u�u�>�3�Ͽ�&����Q��^�Oʗ����_�w�}����Ӏ��`#��t:����c�a�3�
�e��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���d�e�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��h_�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������V��c1��M���8�b�o����0���s���@��V�����2�7�1�g�c�g�5���<����F�D�����%�&�2�6�2��#���H˹��^9��T��!�����n�u�w�.����Y����Z��S
��F���u����l�}�Wϭ�����T��Q��F܊�e�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����U��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%����K����	F��s1��2������u�d�}�������9F������2�%�3�
�c��F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����3�����:�!�"��@���H�ד�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�1��9���=����A��1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������l_��B1�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����/����U��V��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)��������l ��\�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)��������F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�%�)��������U��G]��U���
���
��	�%���Mӂ��]��G�U���&�2�4�u�:��(���&����lT��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2�����¹��lT��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2�����¹��lT��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2��(���&����@��V�����a�
�f�o���;���:����g)��_����!�u�|�_�w�}����ӕ��l��h�����`�
�f�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��V��C1�*���g�a�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l��{:��:���m�
�;�0�'��E���&����CT�=��*����
����u�@Ϻ�����O��N�����4�u�8�
��(�E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�g�<�3��m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
� �f�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h]�� ��a�%�u�u���8���&����|4� N�����u�|�_�u�w�4��������9��h]�*��o������!���6�����Y��E��u�u�&�2�6�}����K���� U��G]��U���
���
��	�%���Y����G	�UךU���<�;�9�%�g�o�(ށ�&����P��N�&���������W��Y����G	�UךU���<�;�9�!�'�i�(�������l��N��1��������}�D�������V�=N��U���;�9�%��$�1�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u��/��#ݰ�����l��Q����� �g�c�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����@��C��*��� �f�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�����
�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��GV��*���f�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӏ��K+��c\�� ���a�3�
�c��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��X�����
�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�e��h�� ��c�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����e9��hZ�*��o������!���6�����Y��E��u�u�&�2�6�}����&˹��lR��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-�D�������U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�4����&����CT�=��*����
����u�W������]ǻN�����9�'�!�<�1��Dف�J����g"��x)��*�����}�a�3�*����P���F��P ��U���
�
�
�
�"�i�C���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�<�3��k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�
�
� �c�o����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*ۊ�
�4�!�6�$����I����	F��s1��2������u�f�}�������9F������&�9�!�%�>�;�(��&���5��h"��<������}�c�9� ���Y����F�D�����
�0� �!�$�;�(��&���5��h"��<������}�`�9� ���Y����F�D������-� ��9�(�(�������C9��1��*��
�g�o����0���/����aF� N�����u�|�_�u�w�4��������l ��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����P��N�&���������W������\F��d��Uʦ�2�4�u�8��d����H����\��c*��:���
�����}�������9F������!�%�g�3��o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
� �`�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[�����f�
�f�o���;���:����g)��Y�����:�e�n�u�w�.����Y����S��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��Z�����u��
����2���+������Y��E��u�u�&�2�6�}�(�������9��h[�*���o������!���6���F��@ ��U���_�u�u�<�9�1����4����])��hX�����%�,�0�3��j�(��Cӵ��l*��~-��0����}�a�1� �)�W���s���@��V�����8�
� �`�g�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����3�
�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���`�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӏ��K+��c\�� ���`�3�
�c��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1��9����!�d�m�1��G߁�I����g"��x)��*�����}�u�8�3���B�����Y�����9�
�g�3��m�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�d�3�
�f��C��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��[��#��
� �c�d�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��ي�
� �c�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_��*���
� �c�d�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V��Dي� �c�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����_	��a1�*���c�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӊ��l0��1��*���
�d�o����0���/����aF�N�����u�|�_�u�w�4��������l��^1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������Z9��h�� ��b�%�u�u���8���&����|4�N�����u�|�_�u�w�4����	����9��h��C���%�u�u����>���<����N��
�����e�n�u�u�$�:��������S��B1�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����/����U��]��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)����ǹ��U��Y��G��������4���Y����\��XN�N���u�&�2�4�w�0�(ށ�&�Փ�l �� ^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�3����H����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�;�#�5�F���&����CT�=��*����
����u�W������]ǻN�����9�;�!�=�e�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʻ�!�=�g�3��n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
� �b�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[�����a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����_��B1�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��T��!�����
����_�������V�=N��U���;�9�;�!�?�n����Oʹ��\��c*��:���
�����}�������9F������;�!�=�f�1��A܁�K����g"��x)��*�����}�u�8�3���B�����Y�����c�
� �b�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��F���
�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��]��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�b���������l ��Y�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����A��h�� ��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Bہ�����R��h��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��Y��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���H˹��W��E	��*���m�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lP��Q��M݊�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����9��Q��Gӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����
9��Q��Fߊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����9��Y�����a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����_��B1�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��B1�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Lƹ��l^��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��F���&����CT�=��*����
����u�W������]ǻN�����9�3�
���	����IŹ��l^��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�4����&����T��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������
V��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�2����&����l_��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�$�1����I����F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����H����lR��B1�C���u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������lW��h]�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G��1�����f�
�f�o���;���:����g)��]����!�u�|�_�w�}����ӕ��l��^��*���l�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�_9��G[�����
�a�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��{+��:���`�
� �l�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��d1��1��� �
�g�!��3�(���@�ԓ�F��d:��9�������w�n�W������]ǻN�����9�!�%�b��(�N���	����`2��{!��6�����u�b�3�*����P���F��P ��U���
�d�3�
�o��F��*����|!��h8��!���}�g�1�"�#�}�^�ԜY�ƿ�T�� �����
� �l�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������[��*���l�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lQ��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�&����P��h=����
�&�
�l�m��3���>����F�D�����%�&�2�7�3�k�C��;����r(��N�����4�u�
�4�e�l�(���H����CW�=��*����
����u�FϺ�����O��N�����4�u�:�
��j����I�ѓ�F��d:��9�������w�j��������l�N�����u�:�
�
�o�;�(��N����	F��s1��2������u�e�}�������9F������!�%�f�<�>����JĹ��\��c*��:���
�����}�������9F������!�%�<�<��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʧ�!�<�
� �f�i�(��Cӵ��l*��~-��0����}�a�1� �)�W���s���@��V�����
�
�d�3��m�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�<�
�"�l�@܁�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�g�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
�g�
�6�)����&����S��G]��U���
���
��	�%���Mӂ��]��G�U���&�2�4�u�2�����K����V��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�����&�ғ�F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���5�Ԣ�F��1��*���
�
�
� �f�m�(��Cӵ��l*��~-��0����}�b�1� �)�W���s���@��V�����a�3�
�d�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@���
�d�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}����I����W��h�Oʆ�������8���Nӂ��]��G�U���&�2�4�u�:��B���&����l��N��1��������}�@Ϻ�����O��N�����4�u�
�a�b�l����H�ӓ� F��d:��9�������w�o�W������]ǻN�����9�!�%�a��(�F��&���5��h"��<������}�g�9� ���Y����F�D�����
�0� �!�d����O¹��\��c*��:���
�����l��������l�N�����u��-� ��3����K����U��G�� ��m�
�f�o���;���:����g)��_����!�u�|�_�w�}����ӕ��l��1��*��b�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��Q��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��h_�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����4����])��hX�����d�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l5��r-�� ���a�g�3�
�e�o����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����g��!�a��(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�l�G���Y�Ɵ�w9��p'�����u�<�;�9�0�-����M����P	��T��!�����
����_�������V�=N��U���;�9�!�%�a����A����\��N��1��������}�CϺ�����O��N�����4�u�8�
�o�;�(��&����W�=��*����
����u�W������]ǻN�����9�!�%�b��(�F�������VF��d:��9�������w�i��������l�N�����u�%�'�!�%��(�������g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����9�4�
�0�"�3�F�������`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����4�u�%�'�#�/�(݁����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�4�
�2�(����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�%������Y����)��t1��6���u�d�u�:�9�2�G��s���P	��X ��ʸ�a�c��m������J���� T��h]��F���9�
�&�u��}�WϹ�����NǻN��U����o�����}���Y���}3��d:��0������]�}�W���Y����l1��c&��U�����n�u�w�}�WϺ�¹��w2��N��!����_�u�u�w�}����.����\��y:��0���n�u�u�%�%�}�}���Y���P
��N��U���
���n�w�}�W�������\��yN��1�����_�u�w�}�W���I����}F��s1��2������u�d�}�������9F�N��U���d�o��u���8���&����|4�_�����:�e�n�u�w�}�WϽ�Y�ƅ�5��h"��<��u�u�u�u�3�(�W���,�Ɵ�w9��p'��#����u�f�u�8�3���Y��ƹF��Y
�����;�;�n�_�w�}����������X��Fҳ�e�3� �
�e�.�Dݰ�&�ԓ�l��h
��U���u�u�2�;�%�>�_���Y���/��N��!����_�u�u�w�}�"���-����	F��c+��'�ߊu�u�u�u�>�m� ���1����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�:�!����Mϗ�-����O��N�����u�_�u�u�w�}���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N����o��u����>���<����N��
�����e�n�u�u�w�}����Y�ƃ�gF��s1��2������u�d�}�������]ǻN�����:�%�;�;�l�W�W�������]����E���f�3�e�3�:��E���J����9��~=ךU���0�0�<�u�]�}�W���Y���/��r)��N���u�u�u����6���Cӯ��v!��d��U���u�1�;�
��	�W���7����a]ǻN��U���<�d����g�>���>����F�N�����
���u�w��2���Y��ƹF��X��]���u�u�u�1�9�}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��Y_��U���������4���Y����W	��C��\�ߊu�u�u�u�'�2���0�Ɵ�w9��p'��#����u�a�1� �)�W���s���F�S��U��� �u��
���(���-���F��@ ��U���|�_�u�u�9�}��������9lǑU�����u�3�e�3�3��E���J���� T��h�����%� �u�u�8�-����Y����_����*���1�f�;�
�e�.�D݁�&����l��=N��U���0�<�u�4�w�W�W���Y�ƅ�[�BךU���u�u� �
���W���J���F�N��ڊ���u�k�d�q�W���Y����Z��`'��=��u�g�_�u�w�}�W�������g.�	N�\���u�%�'�u�6�}�}���Y���P
��
P�����>�_�u�u�w�}����Y����C9��CBךU���u�u�<�e�j�}��������l��=N��U���u�<�d�h�w�/�(���H�֓�JǻN��U���0�h�u�'��(�F�����ƹF�N�����h�u�'�
�"�l�G���P��ƹF��h^�����f�;�
�g�$�n�(ށ�����C9��T�����;�;�u��g�d�D׸�I����_9��Y��G���f�
�
�4��.�}���Y����A��Z��]���u�u�u��w�c�F�ԜY���F��z1��4���h�u�y�u�w�}�WϺ�ù��w2��
P��G�ߊu�u�u�u�>�l� ���1��� T�N��U���1� �
���}�I��P�����CN�����u�u�u�u�3�3�W�������F9��1��Y���u�u�u�1�9�}�IϹ�	����U��G_�U���u�u�1� �w�c��������9��UװU���3�e�3�8��o�������9��T�����;�;�u��g�d�D׸�I����C9��Y��G���d�d�u�u�0�3�������9F�N��U���h�u�y�u�w�}�Wϐ�4����t#�	N����u�u�u�<�g�
�3���D����l�N��Uʱ�;�
���w�c�D��Y���F��X��"����h�u�|�w�}����Y����l�N��Uʱ�;�u�k�2�'�;�(��&����F�N�����u�k�2�%�1��C݁�H���F�N�����u�k�2�%�1��C݁�	����l�N��Uʱ� �u�k�2�'�;�(��&���9l�N��E���8�
�g�&�d�3�(ށ�&�����G������e�l�f�1�m����&�Ԣ�lU��D1��D���u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���|�u�u�%�%�}����s���F�S��U��'�2�d�c�]�}�W���Y����[�^ ��9���;�0�l�0�f�W�W���Y�ƣ�P	��S����c�
� �d�o�2����U���F�
����u�8�
�`�1��Cׁ�K��ƓF�Q1�����
�g�&�f�9��(ށ�N����\��Y��U���e�l�f�3�g�;����K������1�U���2�;�'�6�:�-�_���Y���/��
P��Y���u�u�u����6���D����9F�N��U���e����j�}�E�ԜY���F��Y_��<���u�k�f�y�w�}�W�������d/��N��U���u�u�%�'�w�<�W�ԜY���F��Y^��Kʧ�2�d�c�_�w�}�W������F��h>�����0�l�0�e�]�}�W���Y����W�	N����
� �d�f�8�>���Y���F��X��H���8�
�m�3��h�(��B���F��1�����g�&�f�;���(��CӅ��C	��Y��3��l�f�3�e�1�0�(���
����@9��d��Uʲ�;�'�6�8�'�u�W���Y����wF�_�U���u�u�����2��Y��ƹF�N��������h�w�o�}���Y���W��h9��!���k�f�y�u�w�}�WϺ�����w2��
P��\���u�%�'�u�6�}�}���Y���W��S����d�c�_�u�w�}�W���H���Z��{"�����l�0�d�_�w�}�W���	����[�C��B؊� �d�m�:�4�9�[���Y�����CN��U���
�g�3�
�b��E��s��ƓF�C����� �'�;�u�#�)�Wǿ�&����@�X�����!�!�u�4�?�3�Y��s���R��d1�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�4������E�ƭ�l5��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�u�w�}�W���Y���F�N�����
�&�u�h�6��$������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u�'�/����&ù��V��D��ʥ�:�0�&�u�z�}�WϿ�&����A��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�4��8����I����TF������!�9�f�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����֓�@��G��U���;�_�u�u�w�}�W���Y���F��h�� ���e�%�0�u�j�;�(���<����G9��h\�� ��e�
�f�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����!�'�
�
�%�:�����Ƽ�\��D@��X���u�4�
�0�"�3�F�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��*��� �;�d�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�e�1�0�F���PӒ��]FǻN��U���u�u�u�u�w�}��������9��R	��Hʧ�2�d�d�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����!�'�
�
�%�:�����Ƽ�\��D@��X���u�4�
�0�"�3�E�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��*��� �;�g�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�e�1�0�F���PӒ��]FǻN��U���u�u�u�u�w�}��������9��R	��Hʧ�2�d�`�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����!�'�
�
�%�:�����Ƽ�\��D@��X���u�4�
�0�"�3�D�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��*��� �;�f�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�e�1�0�F���PӒ��]FǻN��U���u�u�u�u�w�}�������� 9��R	��Hʳ�
���g��)�A݁�&����_��G]�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����T��E�����x�_�u�u�%�>��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�r�p�}����Y���F�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��k�^�����ƹF�N��U���u�u�:�9�/�	�8���M˹��T9��[��Hʷ�:�
��,�"��O���&����l��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��P�Ƹ�VǻN��U���u�u�u�u�;��9�������^��h\�����f�m�i�u�;��9�������^��h\�� ��g�%�n�u�w�}�W���Y�����q+��7���:�!� �
�`�m���E�ƪ�l5��r-�� ���e�
�
� �n�k���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�0�u�;�w�2�_ǿ�&����GF�V�����
�:�<�
�~�t�W������F�N��U���u�9������������lV��h_��Hʼ�
�$�f�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��hZ��\ʡ�0�_�u�u�w�}�W���Y�ƪ�l5��r-�� ���a�
�0�
�e�m�K���*����v%��B��AҊ� �c�e�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��F���;�u�:�}�>�����&ǹ��R��R�����g�%�u�u�'�>�����ד�O������u�u�u�u�w�}�Wϸ�&����gT��B��@���'�2�d�c�w�`����4����])��hX��G���
�m�
�f�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��D��\���!�0�_�u�w�}�W���Y���U5��z;��G���!�m�
�
�2��E��E�ƪ�l��{:��:���m�
�
� �d�k���Y���F�N��U���8�
�f�'�0�l�A���DӒ��lS��Q��Eڊ�g�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǻN��Xʴ�&�2�u�'�4�.�Y��s���C��R��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������A�C�����u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���H����^9��G�����_�u�u�u�w�}�W���Y����~3��N!��*���!�%�,�f��8�(��L���T��Q��F܊�g�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǻN��Xʴ�&�2�u�'�4�.�Y��s���C��R��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������A�C�����u�u�u�u�w�;�_�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9��N��U���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���b�3�8�c�~�t����s���F�N��U���'�2�d�`�k�}��������l��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y�����T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��F���|�!�0�_�w�}�W���Y���F��P1�D��u�'�
� �f�k���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�l�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����S�G�����u�u�u�u�w�}�W�������P�
N�����
�f�
�g�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�!�0�_�w�}�W���Y���F��[1�����<�'�2�d�g�}�Jϭ�����W��h��M���%�n�u�u�w�}�W���Y����V
��Z�*���0�
�f�e�k�}��������Z9��hV�*��_�u�u�u�w�}�W���Y����G��1�����d�d�u�h�$�1����@����F9��1��N���u�u�u�u�w�}�Wϭ����� Q��h��*��g�i�u�0��0�D؁�&����S��UךU���u�u�u�u�w�}����N����lW��N�U���
�b�3�
�n��E�ԜY���F�N��Uʡ�%�b�
�0��o�O��Y����U��B1�@���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���u�0�!�&�6�8�_���7����^O��QN��ʦ�4�0�8�6�>�8�W��Y����C9��h��*���<�;�%�:�w�}����
����C9��V��U����
�&�y�6���ԜY�Ʈ�T��N��U���6�&�u�%������
���F�N��U���;�4�
��$�l����I���9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_���
����[��G1�����9�2�6�e�~�t����s���F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ۊ�&�
�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GT��D��U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��F���8�g�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӈ��`2��C]�����u�k�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����*����Z�V��!���a�3�8�f�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��ފ�&�
�u�k�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������l ��R������&�`�3�:�i�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�a�;���s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���ځ�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�
�$��W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�@�������F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$���Ź��^9��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�����Y���F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���A����lQ��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���ׁ�
����X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����l ��hV�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$���ʹ��^9��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��1����_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ӊ�&�
�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GW��Q��L��u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�d�n�w�}�W���Y���F��[��U���u�u�u�u�w�}�W�������l ��R������&�d�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:�����3�8�d�u�i�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d��.�(��s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!�e�;���Y���F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���H����^9��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$����Փ�@��N��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�%������DӇ��`2��C_�����d�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�e�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�f�h�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�`�3�:�l�L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���u�u�0�1�>�f�W���Y���F��_������&�d�
�$��C��Y���F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�V��&���8�i�u�%����������]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	���&����S�	NךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�d�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l�� 1����u�k�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�`�W�W���Y���F�N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�`�;���B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�m�3�8�f�}�I�ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$����ޓ�@�� UךU���u�u�u�u�w�}�������F�N��Uʢ�0�u�%���)�N�������X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�
���F�N��U���u�u�u�4������E�ƭ�l5��D�*���
�m�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����V��D��L��u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ۊ�&�
�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�g�
�&��d�}���Y���F�N�����<�n�u�u�w�}�W�������\��E��K���u�u�u�u�w�}�W�������l ��R��W���������/���!��ƹF�N�����4�0�_�u�w�3�W�������9l�N�U���1�;�u�&�>�3�������KǻN�����;�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B�����y�4�
�<��.����&����l ��h_����u�0�<�_�w�}�W������]	�������!�9�2�6�f�`��������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����_�G�����_�u�u�u�w�}�W�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�:�2�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������]F��X�����x�u�u�4��9����
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�|�u�w�?����Y���F��QN�����}�%�6�;�#�1����H����C9��V��\ʴ�1�}�%�6�9�)���������D�����
��&�d�1�0�G���Y����l�N��U���u�4�
�1�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���'�4�,�4�$�:�W�������K��N�����0�1�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��W��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����V��D��L���u�=�;�_�w�}�W���Y�ƭ�l��S��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-���� ���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������G��h^�����;�%�:�0�$�}�Z���YӇ��A��E ��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�o�(���&���U5��r"��!���
�a�g�3��o�E���UӇ��A��E ��*���2�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��E���8�d�|�|�#�8�W���Y���F������'�
�u�h�1��2���-����R��h��D��
�f�_�u�w�}�W������F�N��Uʴ�
�0� �;�g�a�W�������]9��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������@��YN�����&�u�x�u�w�<�(�������l��^	�����u�u�'�6�$�u����UӔ��lW��N��*���
�&�$���)�G���������E�����
�'�2�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���e�3�8�d�~�t����Y���F�N��U���'�!�'�
�w�`����H����F�N�����u�u�u�u�w�}�WϿ�&����A��R�����0� �;�d�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����
�u�&�<�9�-����
���9F������'�
�
�&�>�3����Y�Ƽ�\��DF����`�u�%�6�{�<�(���&����l5��D�*���
�l�u�%�%�)����&����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���I����lW��G�����_�u�u�u�w�}�W�������]9��S�����c�n�u�u�w�}����Y���F�N��U���'�!�'�
�w�`��������lT��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�/����&�ƭ�@�������{�x�_�u�w�-��������R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�e�3�8�f�q����4����])��hX��G���
�d�`�%�{�<�(�������l��PGךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӇ��A��E ��U��3�
���e����&����lW��1��N���u�u�u�0�$�}�W���Y���F��G1�����
�u�h�4��8����J����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�5�9�F������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��^�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�d�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@Ӈ��Z��G�����u�x�u�u�6���������
9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�4�
�:�$��ށ�Y�ƭ�l%��Q��Aʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@Ӈ��Z��G�����u�x�u�u�6���������
9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�4�
�:�$��ށ�Y�ƭ�l%��Q��D���:�;�:�d�~�f�W�������A	��D����u�x�u�%�$�:����H����@��YN�����&�u�x�u�w�<�(���&����Q��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��D��i�u�4�
�8�.�(���&���R��d1����u�:�;�:�f�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����g�i�u�4��2����¹��F��h-�����d�u�:�;�8�l�^��Y����]��E����_�u�u�x�w�-��������
T��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��W�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����d�g�i�u�6�����&����F�V��&���8�d�u�:�9�2�F���B����������n�_�u�u�z�}��������lT�������%�:�0�&�w�p�W�������T9��S1�G���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�g�g�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��Z�����;�%�:�0�$�}�Z���YӇ��@��U
��G���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�g�a�k�}��������_��N������3�8�b�3�*����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��\�����;�%�:�0�$�}�Z���YӇ��@��U
��G���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�g�g�k�}��������_��N������3�8�d�w�2����H���9F���U���6�&�n�_�w�}�Z���	����l��h]����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�f�u�j�u����&����F��@ ��U���h�4�
�:�$��ށ�P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Bފ�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�b�u�j�u��������EW��S�����
�&�}�l�3�*����@����F�R �����0�&�_�_�w�}�ZϿ�&����Q��V�����;�%�:�0�$�}�Z���YӇ��@��U
��CҊ�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�i�w�<�(���
����9��
N��*���3�8�g�1� �)�W���B����������n�_�u�u�z�}��������lQ��V�����'�6�&�{�z�W�W���	����l��hY�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����b�u�h�}�'�>�����ד�[��G1��*���}�u�:�;�8�k�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����������^	�����0�&�u�x�w�}��������W9��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��i�u�4�
�8�.�(���&���R��d1����1�"�!�u�~�f�W�������A	��D����u�x�u�%�$�:����@�ƭ�@�������{�x�_�u�w�-��������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�l�|�]�}�W���Y����V��=dךU���x�4�
�<��.����&����l ��hW�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�d�
�&����������PF��G�����4�
�<�
�3��O�ԜY�Ʈ�T��N��U���<�u�4�
�>�����A�Ƹ�V�N��U���u�u�4�
�>�����*����V��D��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��E���8�l�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��.����&����l ��h_����2�u�'�6�$�s�Z�ԜY�ƭ�l��h�����
�!�d�3�:�l�(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��_�����e�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���d�
�&�
�g�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9��\�����d�4�&�2�w�/����W���F�V�����&�$��
�#�o����H¹��@��h����%�:�0�&�6��������� OǻN�����_�u�u�u�w�;�_���
����W�� ]�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�d�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�d��.�(��E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�g�6�.��������@H�d��Uʴ�
�<�
�&�&��(���J����lW��V�����'�6�o�%�8�8�ǿ�&����Q��V����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�d�
�$��E��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�F܁�
����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�d�
�$��DϿ�
����C��R��U���u�u�4�
�>�����*����R��D��F���&�2�
�'�4�g��������C9��P1����g�_�u�u�2�4�}���Y���Z �V�����1�
�l�|�#�8�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
����U��]��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�l�(���&����@��YN�����&�u�x�u�w�<�(���&����l5��D�*���
�`�4�&�0�����CӖ��P�������7�1�d�c�]�}�W������F�N��U´�
�<�
�1��m�^Ϫ���ƹF�N��U���%�&�2�6�2��#���HŹ��^9��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���HĹ��^9�������%�:�0�&�w�p�W�������T9��R��!���d�
�&�
�a�<����&����\��E�����%�&�2�7�3�o�E�ԜY�Ʈ�T��N��U���<�u�4�
�>�����I����[��=N��U���u�u�u�%�$�:����&����GW��Q��D���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GW��Q��D���&�<�;�%�8�8����T�����D�����
��&�d��.�(�������]9��X��U���6�&�}�%�$�:����K���F�U�����u�u�u�<�w�<�(���&����U�����ߊu�u�u�u�w�}��������B9��h��M���8�d�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�m�3�:�l�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��*���
�u�&�<�9�-����
���9F������6�0�
��$�l����I����Z��G��U���'�6�&�}�'�.��������9F����ߊu�u�u�u�1�u��������lU�����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�e�����@����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�e�1�0�F���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ي�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�D����ԓ�@��Y1�����u�'�6�&��-��������OǻN�����_�u�u�u�w�;�_���
����W��G�����_�u�u�u�w�}�W���
����@��d:��ي�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��CZ�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�c�;��������]9��X��U���6�&�}�%�$�:����A��ƹF��R	�����u�u�u�3��-��������O��_�����u�u�u�u�w�-��������`2��CZ�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GS��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�`�3�:�i��������\������}�%�&�2�5�9�F��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:��ߊ�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����l ��hX�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�b�3�8�a�<����&����\��E�����%�&�2�7�3�j�^���Yӄ��ZǻN��U���3�}�%�&�0�?���PӒ��]FǻN��U���u�u�%�&�0�>����-����l ��hX��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��CY�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���A����lQ��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=�����3�8�b�4�$�:�(�������A	��D�����2�7�1�g�c�W�W�������F�N�����4�
�<�
�3��E�������9F�N��U���u�%�&�2�4�8�(���
�ޓ�@��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F��������!�a��(�F��&���F��Z��B���
�e�g�%�w�3�W���&����T��G�U���6�
� ���8���&����U��\��F��u�u�u�u�w�4�(�������l_��h_�����}�0�
�8�d��(���&����V�
N��R���9�0�_�u�w�}�W���&����
9��Q��A܊�f�_�u�u�;��2���:����C��Y��*ۊ�
� �d�l�'�}�J���D͏��A��C1�U���0�&�k�x�~�W�W�������w$��|�����f�
�
�
��(�F���	���l�N��Uʴ�
�:�&�
�!�o�Gϩ�����_9��r*��6���!� �
�b�2�l�F���&����CV�N��R��u�9�0�_�w�}�W�������w$��|�����f�
�
�
�l�}�Wϸ�&����p2��C1�C���3�
�g�
�d�a�W���Y��� ��d+��6���!�d�m�'�0�l�@������@��C��B���'�2�d�g��t�J���^�Ʃ�@�N��U���&�9�!�%�g�4����Kù��l�N��*����� �
�g����O����[�N��U���4�
�:�&��+�E��������h[�����b�
�g�e�w�}�F�������9F�N��U���
�c�n�u�w�;�(���<����G9��1��*��
�e�i�u�g�c����
����F��_��H��r�n�u�u�1��2���-����R��Q��Eڊ�f�i�u�u�w�}�Wϸ�&����gT��B��@���'�2�d�c�w�5����*����v%��B��AҊ� �c�e�%��t�J���^�Ʃ�@�N��U���6�
������������9��UךU��������)�Bہ�&����V��G]��H�ߊu�u�u�u�%����I����D��F������,� �
�o�/���M����[�I�����u�u�u�u�w�/���O���F��h=��0��� �
�m�3��k�(��E���X��h�����y�:�=�'�j�z�P��Y����`9��{+��:���`�
� �l�c�-�W��s���F�V�����
�#�g�e� �8�WǸ�&����p2��C1�*���l�a�%�}�~�`�P���Y����l�N��Uʼ�
�!�!����(��Y����`9��u;��9���'�
�g�3��m�(��E�ƥ�l6��P�����0�d�_�u�w�����H����lU��B1�L���u�h�_�u�w�}�W���)����]��1��Eʢ�0�u�!�%�`����M����O�I�\ʰ�&�u�u�u�w�}����H����F�Q=�����
�e�
�
�"�e�A���Y���F�N������'�;�0�n�8�Fϩ�����^��1����l�}�|�h�p�z�W������F�N����c�_�u�u��%�3�������l��^ �����b�
�d�i�w�8�(��B��� ��O#��!ػ� �
�g�g�1��F���	���l�N��Uʳ�
���g��)�A݁����� 9�������0�
�8�m�1��F���	����[�I�����u�u�u�u�w�>�(���=����A��1��G���2�d�g�n�w�}����4����])��hX�����d�f�%�u�j�-�%�������l ��_�*���_�u�u��/��#ݰ�����l��R��#���3�
�d�d�'�}�Jϭ�����Z��R��¦�2�0�}�%�4�3����H˹��u ��E�����1�%��&�;��C���&����l��UךU����-� ��9�(�(�������g��h��D��
�f�i�u�w�}�W�������l��h�����&�
� �d�b��Dϩ�����V
��Z��؊� �d�b�
�e�m�W���H����_��=N��U���u�0�
�8��o����I�ӓ� ]ǻN��&��� ��;� ��h�E���&����CU�
NךU���u�u��-��	����&�ӓ�F9��1��U���;�}�0�
�:�o����A����V�
N��R���9�0�_�u�w�}�W���>����K��C�����d�n�u�u�1��:���K����lP��Q��C܊�d�i�u�
�2�(���&����R��UךU����-� ��9�(�(�������C9��1��*��
�g�i�u�#�����&����\��Y�����4�
�:�&��+�O��Y�ƹ�@��R
��*��� �!�&�3��e�(��P���F��h��9����!�c�
�9�;�#���&����^��N�U���u�u�u�'�#�l����
����@��B1�E���u�=�;�}�2���������Q��G\��\��r�r�u�9�2�W�W���Y�ƿ�_9��G1�����`�
�f�_�w�}�$���,����|��Z��*���f�c�%�u�j�W�W���Y�ƪ�l��{:��:���m�
� �f�c�-�W����ο�_9��GV��*���f�e�%�}�~�`�P���Y����l�N��Uʼ�
��2�<�$�e���s���U5��z;��G���!�m�
� �d�i����DӖ��V��C1�*���f�g�%�n�w�}����4����])��hV�����-�
�
�
�"�o�E���Y����G��X	��*���!�'�&�2�2�u��������EW��(��3���u�<�;�1�'�����&�ԓ�F9��1��\��u�u�3�
���E�������Z��G:�����
�b�
�f�k�}�W���Y����V��h��*���4�!�6�&��(�E���	�ƻ�V�D�����
�d�3�
�`��E��Y���O��[�����u�u�u�0��0�(�������9��dךU���x�2�%�3��n�(�������]F��X�����x�u�u�2�'�;�(��&����@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q�����ƭ�l��h�����
�!�
�&��q��������V��c1��Dۊ�&�
�e�u�'�.��������l��1����y�4�
�<��.����&����l ��h_�U���&�2�6�0��	���&����P�N�����;�u�u�u�w�4�W�������C9��Y�����6�d�h�4��8�^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�d�
�$��G����έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���:�u�4�
�8�.�(�������F��h��*���$��
�!�d�;���PӉ����T�����2�6�d�h�6�����
����g9��Y�����c�u�'�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����u�u�%�6�9�)�������O��_�����u�u�u�u�w�/�(���H�֓�VF������!�9�2�6�g�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��D߁����R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������F9��1��U���<�;�%�:�2�.�W��Y����A��B1�E���
�&�<�;�'�2�W�������@N��h��*���$��
�!��.�(������W�E��D��u�9������������l��h_�� ��l�%�y�4��4�(�������@��Q��A����-� ���)�:������� _��R	��F���u�%�&�2�4�8�(���
����U��]����<�
�&�$���ׁ�
������D�����
��&�d��.�(��s���Q��Yd��U���u�<�u�}�'�>��������lW������6�0�
��$�l�(���&�����YNךU���u�u�u�u�%����I����[��R	��B��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������F9��1��U��3�
���.�(�(�������lU��E��D��n�u�u�u�w�8����Q�έ�l��D�����
�u�u�%�$�:����&����GS��D��\ʺ�u�4�
�:�$�����&���R��^	������
�!�
�$��^�������9F�N��U���u�'�
� �f�m����DӔ��lW��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���ށ�
����F��R ��U���u�u�u�u�0�-����Jù��Z�T��0����� �%�#�n�(���&¹��lW��h����u�u�u�9�2�W�W���Y���F��G1��*��
�e�i�u���/���!����k>��o6��-�������l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����A��B1�E���u�&�<�;�'�2����Y��ƹF��E�� ��e�%�
�&�>�3����Y�Ƽ�\��DF��*���
�&�$���)�(���&����]9��h]����d�`�u����4�������l ��^�����4�
�<�
�$�,�$���ƹ��^9����&�����!�`��(�N���	����C9��P1������&�d�
�$��D���	����l��F1��*���
�&�
�y�6�����
����g9��V�����b�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��DҊ�&�
�b�|�#�8�W���Y���F�	��*���d�e�%�u�j�<�(���
���� T��^�E��_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����U��^��D��u��������&����R��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�/�(���H�֓�F���*��n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W�������F9��1��U��3�
����(�(��&����V��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�/�(���H�֓�F���#���n�u�u�u�w�8����Y���F�N����� �d�e�%�w�`�U���!����k>��o6��-���������U�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�P�����f�
�e�4�$�:�W�������K��N�����3�
�f�
�g�<����&����\��E�����;��
�y�6�����
����g9�� 1����u�%�&�2�4�8�(���
�ғ�@��N��*����g��!�o��(���&����F��h,��1���0�8�g�
������J���R��^	������
�!�f�1�0�F���Y����V��=N��U���u�3�}�4��2��������F�V�����&�$��
�#�n����H���G��d��U���u�u�u�2�'�;�(��&���F��h,��1���0�8�g�
������J����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�2�%�3��n�(��E�ƥ�l0��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�/�(���H�Г�F�������;� �
�c�o����H����9F�N��U���0�_�u�u�w�}�W�������lW��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������9�������%�:�0�&�w�p�W�������F9��1��*���<�;�%�:�w�}����
�Υ�l6��P�����0�e�u�;�3��[Ϭ�����F��h��*���$��
�!��.�(������T9��R��!���a�3�8�f�w�-��������`2��C_�����d�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N�����
�f�
�d�k�}����&��ƹF�N�����u�}�%�6�9�)���������D�����
��&�b�1�0�A�������9F�N��U���u�'�
� �f�k����Dӏ��c*��V��*Ҋ�
�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��F���!�0�u�u�w�}�W���YӁ��l ��]�����h�'�2�d�b�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��Dف�H���>��o6��-���������/���!����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�'�
� �f�o�����ƭ�@�������{�x�_�u�w�/�(���H�ԓ�C��R1�����
�'�6�o�'�2��������T9��R��!���d�
�&�
�g�}����J����lW��B�����8�d�
�
�2��D��Y����G��1�����d�d�y�&�;�)��������lW��B�����8�f�
�
�2��D��Y����Z��D��&���!�g�3�8�f�q��������V��c1��D݊�&�
�c�_�w�}����s���F�^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�a�t����Y���F�N��U���
� �d�g�8�>����DӇ��P	��C1��@��_�u�u�u�w�1����Qۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���;�u�4�
�8�.�(���&���@��C��L���'�2�d�d�~�<����	����@��A_��U���0�
�8�f������J���R��Y��]���6�;�!�9�f�m�Jϭ�����V��h��*��e�|�|�!�2�}�W���Y���F��E�� ��g�:�6�1�w�`��������_��UךU���u�u�9�<�w�u��������_	��T1�Hʴ�
�<�
�&�&��(���K����lW����U´�
�:�&�
�!��W�������l��h_�M���;�u�4�
�8�.�(���&���@��C��D���'�2�d�e�~�<����	����@��A_��U���0�
�8�g������J���R�������!�9�d�e�j�.����	�ߓ�l��h_�C���;�u�4�
�8�.�(���&���@��C��B���'�2�d�g�~�t����Y���F�N��U���
� �d�g�8�>����DӇ��P	��C1��@��_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����U��\�����0�i�u�%�4�3����L����F�N�����u�u�u�u�w�}�WϹ�	����R��X�����h�w���u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���T��Q��A؊�e�4�&�2�w�/����W���F�P�����a�
�e�4�$�:�(�������A	��D������4�2�
���[Ϸ�&����R��hV��*���'�2�d�c�w�-��������`2��C_�����d�y�!�%�`�����K���@��C��D���'�2�d�e�{�.����	�֓�l��h_�E���0�
�8�g������J���@��C��B���'�2�d�g�{�<�(���&����l5��D�*���
�d�u�%�$�:����&����GW��Q��D���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�c�u�'��<�(���
����T��N�����<�
�&�$����������O��Y
�����:�&�
�#��}�W���&����
9��E��D��|�4�1�}�'�>�����ד�[��R����
�
�0�
�d�o�W���Y������T�����d�e�h�&�;�)��������lW��G��\���=�;�_�u�w�}�W���Y����U��\��E��u�0�
�b�l�}�W���YӃ��Z �F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�6�9�_�������l
��h^��U���
�f�'�2�f�d�^Ͽ��έ�l��D��ۊ�u�u�0�
�:�l�(�������R�V ��]���6�;�!�9�f�m�Jϭ�����V��h��*��e�u�;�u�6�����&����F�D�����l�<�'�2�f�l�^Ͽ��έ�l��D��ۊ�u�u�0�
�:�n�(�������T�N�����u�u�u�u�w�}��������9��R������2�<�&�o�8�F�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�f�t�W������F�N��Uʲ�%�3�
�a��m�K�������A��R1����_�u�u�u�w�1��ԜY���F�N�����
�a�
�e�k�}�/���!����k>��o6��-���������L���Y�������U���u�0�1�%�8�8��Զs���K��E�� ��g�%�u�&�>�3�������KǻN����� �d�g�%��.����	����	F��X��¼�
��'�;�2�d���Y����Z��D��&���!�d�3�8�f�q����N����T9��V����!�%�d�<�%�:�F��Uӕ��l��^��*���
�f�e�u�2����&����T9��X����!�%�b�<�%�:�F��UӇ��@��T��*���&�d�
�&��l�W���
����@��d:�����3�8�d�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�b�3�8�f�t�W������F�N��Uʲ�%�3�
�a��l�K���	����@��A]��F��e�e�n�u�w�}�Wϻ�
���N��h�����:�<�
�u�w�-��������`2��C_�����d�|�4�1��-��������lV���*���'�2�d�l�~�<����	����@��A_��U���0�
�8�d������J���R�������!�9�d�e�j�.����	�֓�l��h_�E���;�u�4�
�8�.�(���&���@��C��L���'�2�d�d�~�<����	����@��A_��U���0�
�8�f������J���F��R ��U���u�u�u�u�0�-����M����Z�V�����
�#�g�e�]�}�W���Y����UF������!�9�2�6�f�`��������V��c1��Dۊ�&�
�e�u�%�u��������_	��T1�Hʴ�
�<�
�&�&��(���K����lW����U´�
�:�&�
�!��W�������CT��^1����d�|�4�1��-��������lV���*���f�
�
�0��n�E����Ƣ�GN��G1�����9�d�e�h�$�1����I����V��_�\���u�=�;�_�w�}�W���Y�ƫ�C9��h_�*��i�u�;���<����&����9F�N��U���0�_�u�u�w�}�W�������lW��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�>�����&ǹ��R��R�����g�%�u�h��`��������J��C����x�|�_�u�w�2�(���I����W��G_��Hʳ�
�� ���8���&����R��F�U���u�:�;�:�g�f�W�������lW��Q��Dۊ�a�i�u�
�6�o�F݁�����l��^�����:�g�|�_�w�}����&�ԓ�F9��1��U��%��9�
�e�;�(��&��� F�N�����u�|�_�u�w�2�(���J����R��GZ��Hʥ��9�
�f�1��C܁�H����W	��C��F��u�u�9�6��l�(���O�ѓ�F������d�
� �c�d�-�_��T����\��XN�N���u�9�6��f����J����[��h8��G��
� �c�l�'�u�GϺ�����U�=N��U���
�
�c�3��d�(��E�Ƽ�e��h_�����b�
�d�g�w�}�W������]ǻN�����
�b�3�
�g�j����DӖ��R
��X�� ��d�
�d�f�w�2����K����F�[��#��
� �d�g��l�K���&����lW��Q��E���%�}�f�x�f�9� ���Y����F�[��#���3�
�g�
�f�a�W����ԓ�l ��^�����f�x�d�1� �)�W���s���_	��a1�����e�
�a�i�w��"���7����V��\�� ��a�%�}�e�3�*����J��ƹF��X��*���a�e�%�u�j�-�!���&����lR��h�F���:�;�:�g�~�W�W�������9��hY�*��i�u�e�u�?�3�_���&����l ��V�����u�%�6�;�#�1�O���PӃ��VF�UךU���:�9�&�
�"�j�D���Y���D��_��]���
�
�f�3��i�(��DӇ��P	��C1��M���|�0�&�u�f�f�W�������@U��B1�F���u�h�w�w� �8�Wǲ�����9��hX�*��h�4�
�:�$��ׁ�?�Ʃ�@�L�U���;�!�=�a�1��N߁�K���V�@��U¡�%�b�
� �n�k����Y����\��h��*���u�9�0�w�u�W�W�������l ��W�����h�w�w�"�2�}����/�ߓ�F9��1��U���%�6�;�!�;�e�1�������W�=N��U���'�&�
� �`�l����D������YN�����
�c�3�
�n��F������]��[�*���0�&�u�e�l�}�Wϰ�����l �� ]�����h�w�w�"�2�}����/����U��Y��D��4�
�:�&��+�D��Y����D��d��Uʻ�!�=�f�3��k�(��E���F��R ������d�
� �a�l����Y����\��h��F��u�9�0�w�u�W�W�������9��hW�*��i�u�d�u�?�3�_���&�ד�F9��1��U���%�6�;�!�;�o�(�������V�=N��U���d�d�d�<�1��Fف�J���9F�N��U���6�;�!�9�e��W����θ�C9��h��F���%�}�|�h�p�z�W������F�N�����d�
� �g�o�-�L���YӖ��V��1��*��
�f�i�u�w�}�W�������]��[�*���=�;�}�8��d����H����V�
N��R���9�0�_�u�w�}�W���&����U��^��D�ߊu�u�
�a�b�l����H�ӓ� F�d��U���u�4�
�:�$�����Iӑ��]F��Z��A���
�d�l�%��t�J���^�Ʃ�@�N��U���9�6��d��(�F��&����F�G1�����
�d�3�
�b��B��Yۖ��R
��D1��*��
�d�f�u�8�3���P����^��1��*��
�f�n�u�w�-�%�������l ��V�����h�}�%�6�9�)���&���_	��a1�����e�
�a�n�w�}����
���� U��B1�G���u�h�}����9�������T��B1�A���}�d�1�"�#�}�F���Y����U��h��F���%�|�_�u�w���������U��W�����h�}�%�6�9�)���&���_	��a1�*���d�d�
�a�l�}�WϮ�+����G9��h��D��
�`�i�u�'��݁�O����V��h�F���:�;�:�f�~�{����MŹ��lW��1��\�ߊu�u�
�0�"�)����&����CU�
N�����;�!�9�d��}�W���&����lR��h�N���u�%��9��o����IĹ��Z�E��D��_�u�u�
�6�o�F܁�����l��S������4�2�
���L���YӖ��R
��Z�� ��l�%�u�h�>��;�������l��d��Uʥ��9�
�c�1��G���	�����u;��9���'�
�m�0�e�/���K��ƹF��h8��G���3�
�e�
�f�a�W���>����K��C�����d�n�u�u�'�4����&����T��N�U���u�u�u�3���2�������9��P1�B���=�;�}�8��n����H����O�I�\ʰ�&�u�u�u�w�}����<����|��^�����b�
�f�_�w�}����&����P��h�����
�e�b�%�w�`�}���Y���R��X ��*���`�`�e�"�2�}����J����9��h_�B���}�|�h�r�p�}����s���F�V�����
�#�`�d�g�W�W�������Z9��D�����3�
�`�
�d�a�W���Y�����T�����d�
�e�u�?�3�_���&����Z9��hZ�*��e�u�u�d�~�8����Y���F��G1�����9�d�
�e�l�}�WϬ��ԓ�l��h�����&�
� �g�o�-�W��s���F�V�����
�#�`�`�g�*��������l��h�� ��m�%�}�|�j�z�P������F�N�����:�&�
�#�b�l�G�ԜY�ƾ�G9��h��D��
�f�i�u�w�}�W�������]��[�*��e�"�0�u�#�-�D���¹��lW�� 1��]���h�r�r�u�;�8�}���Y���R��X ��*���`�a�e�n�w�}��������U��G]��H�ߊu�u�u�u�'�>��������V�������8�
�
�
��(�C���	����[�I�����u�u�u�u�w�<�(���
����S��^����u�0�
�
�����M����[�N��U���4�
�:�&��+�B��I�ƻ�V�C��F���<�<�3�
�e��E��Y���O��[�����u�u�u�%�4�3����Hƹ��V��N�����!�%�d�<�1��F؁�K�����h��M���%�u�'�!�'�h�(�������l��B1�B���|�_�u�u�2����&����G9��hV�*��i�u�&�9�#�-�F�������9����U���6�;�!�9�f�l�L���Yӕ��l��\��*���l�m�%�u�j�W�W���Y�ƪ�l5��r-�� ���a�
�0�
�e�m� ���Yە��l��_��*���
�f�a�e�w�}�F�������9F�N��U���!�%�<�3��m�(��s���@��C��M���1�8�'�4��(�O���	���N��G1�*���b�b�%�u�%�.����	�ד�l ��_�����_�u�u�0��0�Fׁ�&����_��N�U¦�9�!�%�m�>�9��������l^��h����4�
�:�&��+�(���s���@��C��L���3�
�f�
�e�a�WǪ�	����U��Y��Gʭ�'�4�
�:�$��ށ�P���F��[1��ۊ� �`�c�%�w�`�U������� ��O#��!ػ� �
�`�<��-��������9��S�����;�!�9�d��m�^ϻ�
���]ǻN�����8�d�<�
�"�o�C���Y���G��^1�����
�g�
�g�/�/��������_��G�U���&�9�!�%��o����I�Փ�F�F�����<�
� �d�d��EϦ�Ӈ��P	��C1��D��n�u�u�&�;�)�ށ�&����P��N�U¡�%�<�<�3��o�(������C9��Y�����d�n�u�u�$�1����I����F9��1��U��}�0�
�8�f��(���A�ߓ�F��SN�����%�l�<�3��n�(��B�����h��Gۊ�
� �l�a�'�}�J�ԜY���F��h=��0��� �
�a�
�2��E��������h��Gڊ�
�0�
�f�g�m�W���H����_��=N��U���u�0�
�8�f��(���@�ޓ� ]ǻN�����8�g�
�
�"�e�D���Y���G��_�� ��b�%�u�;�w�8�(���H¹��]	��Q��A݊�g�n�u�u�$�1����@����F9��1��U��}�8�
�l�1��Nց�KӇ����h��GҊ�
� �m�f�'�t�}���Y����G��h��@���%�u�h�}�2���������l��X�����8�d�3�
�`��E��Y����V
��Z��ۊ� �g�e�%�w�`�_���&ƹ��Z9��Q��A؊�g�4�1�&�;�)�ށ�H����P��G\����u�0�
�8�e�4�(���H����CT�
N�����
�
�d�3��m�F���Y����@��C��*���3�
�e�f�'�t�}���Y����G��h�� ��g�%�u�h��0�(ځ�&����lR��h����&�9�!�%�����O����l�N�����%�e�<�3��o�(��E��ƹF�N��&������!�f�e����H����D��F�����%�l�<�'�0�l�F���P���A�R��U���u�u�u�&�;�)��������
W��G]�U���&�9�!�%�`�4����Oƹ��Z���*���3�
�m�
�e�<�ϭ�����^��h��M���%�|�_�u�w�8�(���M¹��U��\��F��u�u�u�u�w�<�(���
���� T��q-�E��"�0�u�&�;�)��������lW��F�U���d�|�0�&�w�}�W���YӀ��G��1�G���3�
�l�
�d�W�W�������CS��^1��*��
�f�i�u�w�}�W�������A��^��F���
�m�
�f� �8�Wǭ�����V��h��*��e�e�u�u�f�t����Y���F���*���a�
�
� �n�o���Y����V
��Z�*��� �l�c�%�w�`�}���Y���Z��{"�����l�0�e�"�2�}��������l��R	��F��e�u�u�d�~�8����Y���F��R�����
�
� �l�n�-�L���Yӕ��l��1��*��b�%�u�h�u�� ���Yۀ��K+��c\�� ���g�<�
�%�.�8����I�ӓ� F�V�����
�#�`�a�g�t����Y���9F���*���c�<�3�
�a��E��Y���D��F��*����g��!�o�����-����U�� X��F��4�
�:�&��+�B��I����_��^�����u�0�
�8�`�;�(��J����[�L�����}��-� ��3����K����U��G�� ��m�
�f�h�6�����&����lR��N�����e�n�u�u�$�1����&����lU��h�I���d�u�=�;������-����G9��h�����%�
� �g�a�-�W���	����@��A_��A��u�9�0�w�u�W�W�������C^��B1�Mӊ�g�i�u�&�;�)�ف�����9�������!�%�
� �f�e�(��B�����h��M���3�
�m�
�e�a�Wǭ�����9��Q��CҊ�g�:�u�0��0�@�������9��UךU���0�
�8�
�"�h�G���Y���D��_��]���-� ��;�"��B���&����C��B1�M���u�u�%�6�9�)���&����F��D��E��u�u�&�9�#�-�ށ�����l��S��U���u�u�'�!�>�4����&����CU��_��]���
�
�
�
�"�o�E���Q���A��N�����u�u�u�u�6�����&����lR��d��Uʦ�9�!�%�<��(�F��&���FǻN��U���0�
�d�3��m�D���Y����N��G1��ۊ� �d�f�
�e�m�W���H����_��=N��U���u�%�6�;�#�1�Fځ�I��ƹF��R�����
� �a�m�'�}�J�ԜY���F��C1�����f�
�f�"�2�}��������F9��1��]���h�r�r�u�;�8�}���Y���R��X ��*���`�a�e�_�w�}����&����l��B1�F���u�h�w�w� �8�Wǲ�����9��hX�*��h�4�
�:�$�����I�Ʃ�@�L�U���!�%�d�<�>��(���O�ѓ�F�L�U���;�}�:�
��i����LĹ��[��G1�����9�g�
�|�2�.�W��B�����h_��*���
� �c�d�'�}�J���[ӑ��]F��X��*���3�
�g�
�f�`��������_��h^�����u�d�n�u�w�)��������9��R�����u�u�u�%�4�3����A����D��F�����3�
�e�
�e�m�W���H����_��=N��U���u�%�6�;�#�1�O��s���G��1��*��
�f�i�u�w�}�W�������]��[��3���=�;�}�8�����A����O�I�\ʰ�&�u�u�u�w�}��������_��UךU���8�
�
�
�f�;�(��N����[�L�����}�:�
�
�o�;�(��N����F��h�����#�f�e�u�;�8�U���s���G��1�����
�f�
�g�k�}�F������_	��a1�����g�
�d�h�6�����&����lV�R��U��n�u�u�!�'�n��������T��G\��H���w�"�0�u�;�>�!��&����^��N�����:�&�
�#�d�m�W�������l�N����
� �`�c�'�}�J���[ӑ��]F��^	��³�
���g��)�Aځ�����l0��h��A���%�|�i�&�0�8�_�������l
��1�\ʰ�&�u�e�n�w�}����M����U��Z��G��u�d�u�=�9�u����ۀ��K+��c\�� ���a�<�
�-���(���K�ԓ�O������4�
�:�&��+�O��PӃ��VF�UךU���8�
�f�3��i�(��E����^��1��*��
�f�s�%�g�m�(ށ�����l��d��Uʡ�%�a�
�
�"�n�C���Y���G��\�� ��c�%�u�u��l�F������� W��G]����u�8�
�a�1��F���	���D�������<�;�1�3���;���6����9��h��*���
� �d�e��o�W���������T�����d�
��|�2�.�W��B�����hZ�����d�f�%�u�j��Uϩ�����Z��SF��*����g��!�a�����	����l ��_�*��u�u�<�;�3�<�(���
����^��G�����w�w�_�u�w�0�(�������U��N�U¡�%�b�
� �f�i�(��_Ӗ��W��1��*��`�%�|�_�w�}����@����W��G\��H���8�
�
� �b�m����Ӓ��lR��Q��E܊�g�n�u�u�#�-�C���&����l��S��U���u�u�4�
�8�.�(���&����[����*���3�
�d�b�'�u�^��^���V
��d��U���u�4�
�:�$��ׁ�B�����h[�����f�
�f�i�w�}�W���YӒ��lT��B1�C���u�=�;�}�:��N���&����CT�N��R��u�9�0�_�w�}�W�������l ��]����u�u�!�%�b����I����[�C�����
�l�
�g�8�}����K����F9��1��\�ߊu�u�8�
�e�;�(��&���FǻN��U���8�
�
� �d�i�������G��_�� ��e�%�}�|�j�z�P������F�N�����c�
� �f�e�-�L���YӒ��lS��Q��Eڊ�g�i�u�!�'�n��������T��G\��ʻ�!�=�
� �d�i����s���G��Z�����2�;�<�3��n�(��E����^��h�����
�g�
�g�6�9����H����l��B1�D���|�_�u�u�:��B���&����CT�
N�����f�'�2�d�a�}��������lW��h�N���u�!�%�`��8��������F9��1��U��}�8�
�
�o�4����O¹������*ۊ�
�l�<�3��k�(��B�����h[�����g�
�g�i�w�3����H����T��G\��ʻ�!�=�d�3��l�(��B�����h[�����a�
�g�i�w�3����K����U��G\��ʻ�!�=�g�3��n�(��B�����h[�����'�4�
�
�"�j�N���Y���G��^1��*��� �c�b�%�w�3�W���&¹��ZU��h��B���%�|�_�u�w�0�(�������9��R�������g��#�k�(�������lW��B1�A���}�u�u�u�8�3���B�����h[�����`�
�g�i�w�)���&����Q��N��ʡ�%�`�
� �`�h����s���G��1��ۊ� �d�`�
�e�a�W��Y����N��T1��D݊� �d�d�
�c�`��������_��q(�����u�e�n�u�w�)��������F9��1��U��w�w�"�0�w�1��������9��S�����;�!�9�m��t����Y���9F���*ߊ�
�
�
� �e�o����D������YN�����
�
� �g�o�-�W���	����@��AV��3���9�0�w�w�]�}�W���&�ד�F9�� 1��U��}�8�
�l�1��Bށ�KӇ����h��D���%�|�_�u�w�0�(�������9��R��]���'�&�
� �`�d����ӈ��_��h��B���%�|�_�u�w�0�(�������9��R��]���
�g�3�
�`��EϿ�Ӓ��lS��Q��G݊�g�n�u�u�#�-�Aہ�����l��S��&��� ��;� ��i��������9��h\�*��m�x�d�1� �)�W���s���G��[�� ��m�:�6�1�w�`��������_��UךU���8�
�c�3��e�(��E����^��1��*��
�g�4�1�#�-�Aځ�����l��d��Uʡ�%�c�
� �`�n����D�θ�C9��h��B���%�u�;�u�:��@���&����CT�=N��U���
�m�3�
�b��������R��X ��*���
�n�u�u�#�-�Aց�����l��S�����c�
� �b�d�-�W���Y����^��B1�F���|�_�u�u�:��F���&����CT�
N�����b�'�2�d�n�}��������lW��h�N���u�!�%�b��(�F�������VF������!�9�`�a�]�}�W���&�Փ�F9��1��U��}�8�
�f�1��Oށ�KӇ����hY�����`�
�g�n�w�}����Nǹ��lW��1��U��}�8�
�a�1��F���	�ƣ���hZ�����d�f�%�|�]�}�W���&�ӓ�F9��[��F��u�u�u�u�w�)�������� U��N�����!�%�b�
�"�l�Fց�K���F�G�����_�u�u�u�w�0�(�������W��UךU���8�
�c�3��j�(��E�ƪ�l��s����
�:�<�!�1��@݁�H����W	��C��F��u�u�!�%�`����I����Z� �����
� �l�c�'�}�ϰ�����l ��W�����_�u�u�8��m����H�ד�F�������;� �
�e�4�(���&����U��^�����u�u�u�:�9�2�G��Y����^��1��*��
�d�i�u��%�3�������l��^ �����b�
�d�g�w�}�W������]ǻN����� �m�d�%�w�`�_���&�Г�V��P�����
�b�
�g�8�}����A����\��Y1�����e�
�g�n�w�}��������_��G\��H���w�"�0�u�$�:����*����2��x��Mފ�;�0�%��e�;�(��&���F��P ��]���6�;�!�9�f��2�������V�=N��U���
�
�d�3��m�F���Y���D��_��]���
�
�b�3��m�@���Y�ƭ�l��D��Ҋ�|�0�&�u�g�f�W�������l��^1��*��
�g�i�u�f�}����Q����e9��h��C���%�u�u�%�4�3����A������RN��W�ߊu�u�8�
��i����&����CT�
N��Wʢ�0�u�9�6��l�(���O�Փ�F�V�����
�#�
��w�1����[���F��G1��Ҋ�
� �c�d�'�}�J���[ӑ��]F��X��*���3�
�a�
�c�`��������_��q(�����u�e�n�u�w�)��������T��G\��H���w�"�0�u�;�>�!���&����CR������!�9�m�e�w�1����[���F��G1�����3�
�g�
�e�a�W��Y����N��T1��L���
�e�
�a�j�<�(���
����9�������w�_�u�u�:��(���L�֓�F�L�U���;�}�<�;�3�;�(���5�Ԣ�F��1��*���
�
�
� �c�i����Gӕ��]��V�����
�#�m��~�}����[����V��U����