-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�u� �2�4��������T��_�[���n�_�&�u�2�8��������l��^	��Ĵ�9�_�0�!�#�}�Gݚ�O�Ҋ�lV��h_�����
�
�:�u�$�W�W�������PNǻN��U���u�u�1�<�#�}�W���Y����T��S��C���u�u�u�u�w�}�W������F������u�h�d�n�]�}�W���Y�����h�����u�u�;�0�2�}�J��K���F�d��Uʥ�'�u�_�u�w�}�W�������F�T��ʦ�1�9�2�6�!�>��������W��X����n�_�u�u�w�}�W���Y���F��^ �����:�<�n�_�w�}�W���Y���F�N��U���u�!�
�:�>�����ۂ��W��N�����u�|�_�u�w�}�W�������F�T��ʦ�1�9�2�6�!�>��������W��X����n�_�u�u�w�}�W���Y���F��^ �����:�<�n�_�w�}�W���Y���F�N��U���u�!�
�:�>�����ۂ��W��N�����u�|�_�u�w�}�W������F�N��U���
�:�<�_�w�}�L����Ʃ�G��Nװ���=�!�6� �2�/�ϱ�Y����P��q��*���d�>�'�
��2�W���s����]��V
��E���%�o�&�1�;�:��������R��C��U���;�:�e�n�]�4��������l��T�����:�<�
�0�#�/��������W	��C��\���!�%�u�0��/����
Ӈ��R�N��U���
�<�0�d�w�;��������l��C��]���1�=�d�1� �)�W���Y����]��Z��Oʸ�8�4�'�,�m�}�}���Y���D��^�E��e�e�e�w�w�}�I���I����V��^�E���u�u�k�w�g�m�G��I����V�d��U��h�u�e�e�g�l�G��H����F��
P��E��e�d�e�d�g�m�U���Y���V��^�D��d�e�w�u�w�}�A��Y����V��_�D��e�y�b�h�w�m�G��I����W��L�M��u�e�e�e�f�m�G��I���9F�W��K���e�e�d�d�g�l�G��U����X�^�E��d�e�d�e�u�}�F��Y����W��_�E��e�y�_�u�w�o�J���I����V��_�E��y�d�u�k�u�m�G��I����V��B��A��u�e�e�d�f�l�F��H���9F�_�H���e�e�d�d�f�m�G��[����[�^�E��e�e�e�d�g�q�F���G����V��_�E��e�w�u�u�w�l�W���[����W��^�D��w�u�l�h�w�m�G��H����V��L�G���k�w�e�e�f�l�G��I���l�N�U��w�e�d�e�g�l�F��H���F�L�E��e�e�d�d�f��W��D���V��_�E��e�d�y�_�w�}�C��Y����V��_�E��e�y�g�u�i��G��I����V��_��U��h�u�e�e�g�m�G��I����FǻN��B��u�e�e�e�g�m�G��I���^�	N��E��d�d�d�e�g�m�[��Y���V��_�D��d�e�w�u�w�}�D���G����W��_�D��d�w�u�d�j�}�G��H����W��_�Y��u�k�w�e�f�m�G��H����J�N��F���k�w�e�d�g�l�G��H���U��
P��E��d�d�d�e�g�l�U���L���V��_�D��e�d�d�y�]�}�W��D���V��^�E��d�e�y�f�w�c�U��H����W��^�W���m�h�u�e�g�l�G��I����D�=N��U��h�u�e�e�f�l�G��I����F��S�W��d�d�d�e�f�m�G��M���D��_�D��e�d�e�w�w�}�W��Y���V��^�D��d�d�w�u�d�`�W��H����V��^�E���a�u�k�w�g�m�G��I����V�d��U��u�k�w�e�g�m�G��I����J�N��U��d�e�d�d�f�m�F���Y���F�_�D��d�e�d�d�{�W�W���A���V��^�D��e�e�e�y�c�}�I���I����W��^�E���u�e�h�u�g�l�G��H����V��NךU���d�h�u�e�f�m�F��H����D�\��K���e�e�e�e�g�m�F��U����X�^�D��d�d�e�e�u�}�W���L���D��^�E��d�e�e�w�w�h�J���I����W��_�E��y�`�u�k�u�m�G��H����W��B��U���`�u�k�w�g�m�G��H����V�[�H���e�d�d�e�f�m�F��[����[�^�E��d�d�d�d�f�q�}���Y���F�_�D��e�d�e�d�{�k�W���[����W��_�D��w�u�g�h�w�m�F��H����V��L����u�f�h�u�g�l�G��I����W��N�U��w�e�d�e�g�l�F��I���F�L�D��e�d�d�e�g��W���Y����X�^�E��e�d�d�d�u�}�@��Y����V��^�E��d�y�c�u�i��G��I����W��_��U���u�c�u�k�u�m�F��I����W��B��E��u�e�d�e�g�m�G��H���W�	N��E��d�e�e�e�f�m�[�ԜY����[�^�D��e�e�d�e�g�q�@���G����W��_�D��e�w�u�a�j�}�G��H����W��^�Y�ߊu�u�`�h�w�m�F��I����W��L�B���k�w�e�d�g�l�G��H���Q��
P��E��d�d�e�e�g�m�U���Y���F�L�D��d�d�d�e�f��W��D���W��_�E��d�d�y�m�w�c�U��H����W��_�W���u�u�m�u�i��G��H����V��^��U��h�u�e�d�f�m�F��H����F��S�W��d�d�e�d�g�m�G��s���R�	N��E��d�d�e�d�f�l�[��Y���V��_�D��e�d�w�u�a�`�W��I����V��^�E���_�u�u�b�j�}�G��I����W��^�Y��u�k�w�d�g�m�F��I����J�N��U��e�e�d�e�f�l�F���Y���_��
P��E��e�d�e�d�g�l�U���H���V��^�D��d�e�d�y�n�}�I���H����V��_�D���u�u�u�l�w�c�U��I����V��_�W���a�h�u�e�g�m�G��I����D�[��K���d�e�d�e�f�l�F��U���F��S�W��e�d�d�e�f�l�F��@���D��^�D��e�e�e�w�w�e�J���I����V��_�E��y�_�u�u�n�`�W��I����V��_�D���d�e�h�u�g�m�F��H����V��N�D��u�e�e�d�f�m�G��I���9F�_�U��w�d�e�e�g�l�F��H���U�	N��D��e�d�e�d�f�m�[��M���V��_�E��e�e�e�y�]�}�W��Y���W��_�D��e�e�w�u�g�}�I���H����W��^�E���u�e�u�k�u�l�G��I����V��B��U���d�m�h�u�g�m�F��H����V��N�L��u�e�e�d�f�m�G��H���W��
P��E��d�d�d�d�f�l�U���Y���W�	N��D��e�e�e�d�g�m�[��K���V��^�D��d�d�e�y�f�n�J���I����V��^�D��y�_�u�u�f�}�I���H����V��^�E���u�d�u�k�u�l�F��H����V��B��D���k�w�d�d�g�l�G��I���l�N�B��u�e�e�e�g�m�F��H���W��
P��E��e�e�d�e�f�l�U���H���D��_�E��d�e�e�w�w�}�W��I���V��^�D��d�d�e�y�f�l�J���I����W��^�E��y�d�g�h�w�m�G��H����W��L����u�g�u�k�u�l�F��H����V��B��G���k�w�d�d�g�m�F��I���W��S�W��d�e�e�d�f�l�G��s���T��
P��E��d�e�e�d�g�m�U���K���D��_�E��d�e�e�w�w�o�W���[����V��^�E��w�u�u�u�f�d�J���I����W��^�E��y�d�e�h�w�m�G��H����W��L�D��h�u�e�e�f�m�G��H����FǻN��F���k�w�d�d�f�m�G��H���W��S�W��d�d�d�e�f�l�G��H���F�^�D��d�e�e�e�{�W�W���J���D��_�D��e�e�e�w�w�n�W���[����W��_�E��w�u�f�u�i��F��H����W��^��U���u�d�m�h�w�m�G��H����V��L�D��h�u�e�d�g�m�G��H����F��N��U��d�e�e�d�f�l�G���Y���W��S�W��e�e�d�d�g�l�F��H���F�_�E��d�d�e�d�{�l�D��Y����V��^�D��e�y�_�u�w�i�W���[����V��_�E��w�u�a�u�i��F��I����W��_��U��u�k�w�d�g�m�F��I����J�N��D��h�u�e�d�g�m�G��H����F��N��U��d�e�e�d�f�l�G���Y����X�_�E��e�d�e�e�u�}�W���H���F�_�D��d�d�d�e�{�l�F��Y����V��^�D��d�y�d�g�j�}�G��I����V��^�Y�ߊu�u�`�u�i��F��H����V��_��U���u�k�w�d�g�l�F��H����J�[��K���d�e�e�e�g�l�G��U���F��N��U��d�d�e�d�f�m�F���Y����X�_�D��e�e�d�d�u�}�B���G����V��_�E��e�w�u�u�w�l�N��Y����W��_�D��d�y�d�e�j�}�G��H����W��_�Y��d�h�u�e�f�l�F��I����D�=N��U��u�k�w�d�g�m�F��I����J�]��K���d�e�e�d�g�l�G��U����[�^�E��e�e�e�d�g�q�}���Y����X�_�D��d�e�d�d�u�}�A���G����V��^�D��e�w�u�c�w�c�U��I����W��^�W���u�u�d�m�j�}�G��H����V��_�Y��l�h�u�e�f�l�F��H����D�Y�H���e�d�d�d�f�m�G��[��ƹF� _��K���d�e�d�e�f�l�G��U����[�^�E��d�d�d�d�f�q�F��D���W��_�D��e�e�y�_�w�}�@���G����W��^�D��d�w�u�b�w�c�U��H����V��^�W���b�u�k�w�f�l�G��H����W�d��U��b�h�u�e�f�m�G��I����D�Y�H���e�d�e�e�f�m�F��[����
F�L�D��e�d�d�d�f��W���Y����[�^�D��e�d�d�d�f�q�F��D���W��_�E��d�d�y�d�e�`�W��H����V��_�E���_�u�u�m�w�c�U��H����W��_�W���m�u�k�w�f�l�G��I����V�_�U��w�d�d�d�g�m�G��H���F�V�H���e�d�e�e�g�l�G��[����F�L�D��e�d�d�e�f��W��Y���W��_�E��e�e�w�u�w�}�F��D���W��^�D��d�e�y�d�g�`�W��H����W��^�E���d�d�h�u�g�l�G��H����V��NךU���l�u�k�w�f�l�F��H����V�_�U��w�d�d�d�g�m�G��I���
R�	N��D��d�e�d�d�g�l�[�ԜY����F�L�D��d�e�d�e�f��W��Y���W��_�E��d�e�w�u�n�}�I���H����W��_�E���u�u�u�d�o�`�W��H����W��_�D���d�l�h�u�g�l�F��I����V��N�E��u�e�d�d�g�l�G��I���9F�\�U��w�d�d�e�g�l�G��I���T�	N��D��e�d�e�e�g�m�[��J���V��_�D��e�e�e�y�]�}�W��Y���W��^�D��d�d�w�u�g�}�I���H����W��^�E���u�e�u�k�u�l�F��I����W��B��U���g�b�h�u�g�l�F��I����W��N�M��u�e�d�d�f�m�F��I���V��
P��E��d�d�d�d�g�l�U���Y���V�	N��D��e�e�d�e�f�l�[��H���V��_�D��e�d�d�y�e�o�J���I����W��^�D��y�_�u�u�f�}�I���H����W��_�D���u�d�u�k�u�l�F��H����W��B��D���k�w�d�d�g�l�F��I���l�N�C��u�e�d�d�g�m�F��H���W��
P��E��d�e�e�e�f�l�U���H���D��_�E��e�d�e�w�w�}�W��@���V��_�E��d�d�d�y�e�m�J���I����V��_�D��y�g�d�h�w�m�F��I����W��L����u�g�u�k�u�l�F��H����V��B��G���k�w�d�d�f�l�F��I���T��S�W��d�d�d�e�g�m�G��s���T��
P��E��d�e�d�d�g�m�U���K���D��_�E��e�e�d�w�w�o�W���[����W��_�D��w�u�u�u�e�e�J���I����W��^�D��y�g�l�h�w�m�F��H����W��L�G��h�u�e�d�f�l�G��I����FǻN��F���k�w�d�d�f�m�F��H���T��S�W��d�d�e�e�f�l�F��K���F�_�D��e�d�e�e�{�W�W���J���D��_�D��e�e�d�w�w�n�W���[����W��_�E��w�u�f�u�i��F��H����V��^��U���u�g�b�h�w�m�F��H����V��L�G��h�u�e�d�f�l�G��H����F��N��U��d�d�d�e�g�l�F���Y���T��S�W��d�d�d�d�g�m�G��K���F�_�D��d�d�d�d�{�o�E��Y����W��_�E��d�y�_�u�w�i�W���[����W��^�D��w�u�a�u�i��F��H����V��_��U��u�k�w�d�f�l�F��H����J�N��G��h�u�e�d�f�l�F��I����F�� N��U��d�d�d�d�g�l�F���Y����X�_�D��d�e�d�e�u�}�W���K���F�_�D��d�e�e�e�{�o�G��Y����W��_�E��e�y�g�d�j�}�G��H����W��^�Y�ߊu�u�`�u�i��F��H����W��^��U���u�k�w�d�f�l�F��H����J�Z��K���d�d�d�d�f�l�F��U���F��N��U���h�u�e�d�f�l�F��H����F��N��U��d�d�d�d�f�l�F���Y����X�_�D��d�d�d�d�u�}�W���K���F�_�D��d�d�d�e�{�o�F��Y����W��_�D��d�y�g�g�j�}�G��H����W��_�Y�ߊu�u�c�u�i��F��H����V��^��U��u�k�w�d�f�l�F��H����J�[��K���d�d�d�d�f�m�F��U���F��N��U��d�d�d�d�g�m�F���Y����X�_�D��d�d�e�e�u�}�A���G����W��_�D��d�w�u�u�w�o�N��Y����W��_�D��e�y�g�e�j�}�G��H����V��_�Y��d�h�u�e�f�l�F��H����D�=N��U��u�k�w�d�f�l�F��I����J� ]��K���d�d�d�d�f�m�F��U����[�^�D��d�e�d�e�g�q�}���Y����X�_�D��e�d�e�d�u�}�@���G����W��_�E��d�w�u�b�w�c�U��H����W��^�W���u�u�g�m�j�}�G��H����V��_�Y��l�h�u�e�f�l�F��H����D�V�H���e�d�d�d�f�m�F��[��ƹF�_��K���d�d�d�e�f�l�F��U����[�^�D��e�d�e�e�g�q�E��D���W��_�E��d�d�y�_�w�}�O���G����W��^�E��d�w�u�m�w�c�U��H����W��^�W���m�u�k�w�f�l�F��H����V�d��U��b�h�u�e�f�l�G��H����D�V�H���e�d�d�e�f�m�F��[����
F�L�D��e�e�d�e�f��W���Y����[�^�D��d�e�d�e�g�q�E��D���W��^�E��d�d�y�g�e�`�W��H����W��^�E���_�u�u�l�w�c�U��H����V��_�W���l�u�k�w�f�l�F��I����W�\�U��w�d�d�d�g�l�F��I���F�W�H���e�d�d�e�g�l�F��[����F�L�D��d�d�d�d�g��W��Y���W��^�D��e�d�w�u�w�}�E��D���W��_�E��e�e�y�f�g�`�W��H����V��_�D���f�d�h�u�g�l�F��I����W��NךU���e�u�k�w�f�l�G��H����W�]�U��w�d�d�e�g�m�F��H���R�	N��D��e�e�d�d�f�l�[�ԜY����F�L�D��d�e�e�e�f��W��Y���W��^�E��e�d�w�u�g�}�I���H����W��^�E���u�u�u�f�o�`�W��H����W��_�E���f�l�h�u�g�l�F��I����W��N�E��u�e�d�d�g�m�G��H���9F�]�U��w�d�d�e�g�l�G��I���T�	N��D��e�e�e�e�f�l�[��J���V��_�E��e�e�e�y�]�}�W��Y���W��_�D��d�d�w�u�f�}�I���H����W��_�E���u�d�u�k�u�l�F��H����W��B��U���f�b�h�u�g�l�G��I����W��N�M��u�e�d�e�f�l�G��I��� W��
P��E��e�d�d�e�f�l�U���Y���V�	N��D��d�e�d�e�g�m�[��H���V��^�D��d�d�e�y�d�o�J���I����V��_�D��y�_�u�u�e�}�I���H����W��_�D���u�g�u�k�u�l�F��H����W��B��G���k�w�d�d�f�m�G��I���l�N�C��u�e�d�e�g�m�F��I��� T��
P��E��e�e�e�e�f�l�U���K���D��_�D��d�e�d�w�w�}�W��@���V��^�D��d�d�d�y�d�m�J���I����W��^�E��y�f�d�h�w�m�F��H����W��L����u�f�u�k�u�l�F��I����W��B��F���k�w�d�d�g�l�F��I���U��S�W��d�e�d�e�f�l�G��s��� U��
P��E��e�e�e�e�g�m�U���J���D��_�E��d�e�d�w�w�n�W���[����V��^�E��w�u�u�u�d�e�J���I����V��_�E��y�f�l�h�w�m�F��H����V��L�F��h�u�e�d�f�l�G��H����FǻN��A���k�w�d�e�f�m�F��I���U��S�W��e�d�e�e�f�l�F��J���F�_�D��e�d�e�d�{�W�W���M���D��^�E��e�d�d�w�w�i�W���[����W��_�E��w�u�a�u�i��F��H����W��_��U���u�f�b�h�w�m�F��I����W��L�F��h�u�e�d�f�m�G��I����F��N��U��d�d�d�d�f�l�G���Y���U��S�W��e�e�d�d�g�m�F��J���F�_�E��d�d�d�d�{�n�E��Y����W��^�E��e�y�_�u�w�h�W���[����V��_�D��w�u�`�u�i��F��I����V��^��U���u�k�w�d�g�m�F��H����J�N��F��h�u�e�d�f�m�F��I����F�� N��U��d�d�e�e�f�m�F���Y����X�_�E��d�d�d�e�u�}�W���J���F�_�D��d�e�d�d�{�n�G��Y����V��_�D��e�y�f�d�j�}�G��I����V��_�Y�ߊu�u�c�u�i��F��H����W��^��U��u�k�w�d�g�l�F��I����J�Z��K���d�e�d�e�f�m�G��U���F��N��U��d�e�e�e�f�l�G���Y����X�_�E��d�d�d�d�u�}�A���G����V��_�D��e�w�u�u�w�n�O��Y����V��_�D��e�y�f�l�j�}�G��I����W��_�Y��e�h�u�e�f�m�G��H����D�=N��U��u�k�w�d�g�m�F��I����J� \��K���d�e�e�e�f�m�F��U����[�^�E��e�d�e�e�g�q�}���Y����X�_�D��d�d�e�e�u�}�@���G����W��_�E��d�w�u�b�w�c�U��H����W��_�W���u�u�f�b�j�}�G��H����V��^�Y��m�h�u�e�g�l�G��I����D�Y�H���e�e�d�e�g�l�F��[��ƹF�^��K���d�d�d�e�g�l�F��U����[�^�D��e�e�e�e�f�q�D��D���V��_�E��d�d�y�_�w�}�O���G����W��_�E��e�w�u�m�w�c�U��H����V��^�W���m�u�k�w�f�l�G��H����V�d��U��c�h�u�e�g�l�G��H����D�V�H���e�e�d�e�f�m�G��[����F�L�E��e�e�e�e�f��W���Y����[�^�D��d�e�d�e�f�q�D��D���V��_�E��d�e�y�f�f�`�W��I����W��_�E���_�u�u�l�w�c�U��H����W��_�W���l�u�k�w�f�l�F��H����V�]�U��w�d�d�d�g�l�G��I���F�W�H���e�e�e�e�g�l�G��[����F�L�E��d�d�e�d�f��W��Y���W��^�E��e�d�w�u�w�}�D��D���V��_�D��e�d�y�f�n�`�W��I����W��_�D���a�e�h�u�g�m�G��I����V��NךU���e�u�k�w�f�l�G��I����V�Z�U��w�d�e�d�f�l�F��H���U�	N��D��d�d�d�d�f�m�[�ԜY����F�L�E��d�d�e�e�g��W��Y���W��_�E��e�e�w�u�g�}�I���H����W��^�E���u�u�u�a�`�`�W��I����W��^�D���a�m�h�u�g�m�F��I����V��N�L��u�e�e�d�f�l�G��H���9F�Z�U��w�d�e�e�g�l�F��H���W�	N��D��e�e�d�d�g�m�[��K���V��_�D��d�d�e�y�]�}�W��Y���W��^�E��d�d�w�u�f�}�I���H����V��^�D���u�d�u�k�u�l�G��H����W��B��U���a�c�h�u�g�m�G��I����V��N�B��u�e�e�e�f�m�F��I���W��
P��E��e�e�d�e�f�m�U���Y���_�	N��D��d�d�e�e�f�m�[��I���V��^�E��d�e�d�y�c�l�J���I����W��^�E��y�_�u�u�e�}�I���H����W��^�D���u�g�u�k�u�l�G��I����V��B��G���k�w�d�e�g�l�F��H���l�N�@��u�e�e�e�g�m�F��I���T��
P��E��e�e�e�d�g�m�U���K���D��_�D��e�e�d�w�w�}�W��A���V��_�D��d�d�d�y�c�d�J���I����W��_�E��y�a�e�h�w�m�F��I����W��L����u�f�u�k�u�m�F��H����V��B��F���k�w�e�d�f�m�F��H���R��S�W��d�e�d�e�g�l�F��s���U��
P��E��d�d�d�d�g�l�U���J���D��_�D��e�e�e�w�w�n�W���[����V��^�D��w�u�u�u�c�j�J���I����V��^�E��y�a�m�h�w�m�F��I����V��L�A��h�u�e�d�g�l�G��I����FǻN��A���k�w�e�d�f�m�G��I���R��S�W��d�d�e�e�g�l�G��M���F�_�D��d�e�d�e�{�W�W���M���D��_�E��e�e�d�w�w�i�W���[����V��_�D��w�u�a�u�i��G��I����V��_��U���u�a�c�h�w�m�F��H����W��L�A��h�u�e�d�g�m�F��I����F��N��U��d�e�e�d�f�l�G���Y���R��S�W��d�e�e�d�g�m�G��M���F�_�D��e�e�d�d�{�i�F��Y����W��_�E��e�y�_�u�w�h�W���[����W��^�E��w�u�`�u�i��G��H����W��_��U���u�k�w�e�g�l�G��H����J�N��A���h�u�e�d�f�l�F��H����F��N��U��d�d�d�e�g�l�F���Y����X�^�D��e�d�e�d�u�}�W���M���F�_�E��e�e�d�e�{�i�N��Y����W��_�E��d�y�a�e�j�}�G��H����W��_�Y�ߊu�u�c�u�i��G��H����V��^��U��u�k�w�e�g�l�G��I����J�]��K���e�e�d�d�f�m�G��U���F��N��U��d�e�e�e�f�l�G���Y����X�^�E��e�d�e�d�u�}�A���G����V��_�D��d�w�u�u�w�i�@��Y����V��_�E��d�y�a�m�j�}�G��I����W��^�Y��l�h�u�e�f�m�G��H����D�=N��U��u�k�w�e�g�m�G��H����J� _��K���e�d�d�d�f�l�F��U����[�^�D��d�e�d�e�g�q�}���Y����X�^�D��e�e�e�d�u�}�@���G����W��_�E��d�w�u�b�w�c�U��H����W��^�W���u�u�a�c�j�}�G��H����V��^�Y��b�h�u�e�g�l�F��I����D�Y�H���e�e�d�d�f�m�G��[��ƹF� W��K���e�d�e�d�g�l�F��U����[�^�D��e�d�d�e�f�q�C��D���V��^�E��e�d�y�_�w�}�O���G����W��_�D��d�w�u�m�w�c�U��H����V��^�W���m�u�k�w�g�l�F��H����V�d��U��`�h�u�e�g�m�G��I����D�V�H���e�e�e�e�g�m�G��[����F�L�E��d�d�e�d�f��W���Y����[�^�D��e�d�e�e�g�q�C��D���V��_�E��e�d�y�a�g�`�W��I����V��_�E���_�u�u�l�w�c�U��H����W��^�W���l�u�k�w�g�m�F��I����W�Z�U��w�e�e�d�g�l�G��I���F�W�H���e�e�d�d�g�m�F��[����F�L�E��e�e�e�e�g��W��Y���V��_�D��d�e�w�u�w�}�C��D���V��_�D��d�e�y�a�o�`�W��I����W��_�D���a�l�h�u�g�m�F��I����W��NךU���e�u�k�w�g�m�G��H����W�[�U��w�e�e�e�g�m�G��I���T�	N��E��d�d�d�d�g�l�[�ԜY���� F�L�E��d�e�e�e�g��W��Y���V��_�E��d�e�w�u�g�}�I���I����W��_�D���u�u�u�`�a�`�W��I����W��^�E���`�b�h�u�g�m�G��H����V��N�M��u�e�e�e�f�m�F��I���9F�[�U��w�e�e�e�g�l�F��H���V�	N��E��e�d�e�d�g�m�[��H���V��^�E��e�e�d�y�]�}�W��Y���V��^�E��e�e�w�u�f�}�I���H����W��_�D���u�d�u�k�u�l�F��I����W��B��U���`�`�h�u�f�l�F��H����V��N�C��u�d�d�d�g�l�G��I���W��
P��D��d�e�e�e�g�l�U���Y���^�	N��D��e�d�d�e�g�m�[��@���W��_�E��e�e�d�y�b�m�J���H����V��_�E��y�_�u�u�e�}�I���H����V��^�D���u�g�u�k�u�l�F��I����W��B��G���k�w�d�d�f�l�F��H���l�N�A��u�d�d�e�f�l�G��I���T��
P��D��e�e�d�e�f�m�U���K���D��_�E��e�e�e�w�w�}�W��N���W��^�E��d�d�e�y�b�e�J���H����W��_�D��y�`�l�h�w�l�F��H����W��L����u�f�u�k�u�l�F��H����W��B��F���k�w�d�d�g�l�G��H���S��S�W��d�e�e�d�f�l�F��s���U��
P��D��d�d�d�e�f�m�U���J���D��^�D��e�e�d�w�w�n�W���[����W��_�D��w�u�u�u�b�k�J���H����V��_�E��y�`�b�h�w�l�F��I����V��L�@��h�u�d�d�f�l�F��H����FǻN��F���k�w�d�e�g�m�F��H���S��S�W��e�e�e�e�f�l�G��L���F�_�E��d�d�e�e�{�W�W���M���D��^�E��e�e�d�w�w�i�W���[����W��_�D��w�u�a�u�i��F��H����V��_��U���u�`�`�h�w�l�F��H����V��L�@��h�u�d�d�g�m�G��H����F�� N��U��d�e�e�d�f�l�G���Y���S��S�W��e�e�d�d�f�l�G��L���F�_�E��e�d�e�e�{�h�G��Y����V��^�E��d�y�_�u�w�h�W���[����V��^�D��w�u�`�u�i��F��I����V��^��U���u�k�w�d�g�m�G��I����J�N��@��h�u�d�e�f�l�G��I����F��N��U��e�d�d�d�g�l�F���Y����X�_�D��d�e�d�e�u�}�W���L���F�^�D��e�d�e�d�{�h�O��Y����W��^�D��d�y�`�l�j�}�F��H����V��^�Y�ߊu�u�c�u�i��F��I����W��^��U��u�k�w�d�f�m�G��H����J�\��K���d�d�e�d�f�l�G��U���F��N��U��e�d�e�d�g�l�G���Y����X�_�E��d�e�d�e�u�}�A���G����W��_�E��d�w�u�u�w�h�A��Y����V��^�D��e�y�`�b�j�}�F��I����V��_�Y���m�h�u�d�g�m�G��H����D�=N��U��u�k�w�d�f�l�G��I����J� ^��K���d�d�e�d�f�m�F��U����[�_�D��e�e�e�e�f�q�}���Y����X�_�E��d�d�d�d�u�}�@���G����W��_�D��e�w�u�b�w�c�U��H����W��^�W���u�u�`�`�j�}�F��H����W��_�Y���c�h�u�d�g�l�F��I����D�Y�H���d�e�d�d�g�m�F��[��ƹF� V��K���d�e�d�d�g�l�G��U����[�_�E��e�d�d�e�f�q�B��D���V��^�E��e�d�y�_�w�}�O���G����V��_�D��e�w�u�m�w�c�U��I����V��^�W���m�u�k�w�f�m�G��H����V�d��U���a�h�u�d�g�l�G��I����D�V�H���d�e�d�e�f�m�G��[����F�L�E��d�d�e�d�f��W���Y����[�_�E��d�e�e�d�f�q�B��D���V��_�D��e�d�y�`�n�`�W��I����W��^�E���_�u�u�l�w�c�U��I����V��_�W���l�u�k�w�f�m�F��H����W�[�U��w�d�e�e�f�m�G��H���F�W�H���d�e�e�d�f�l�F��[����F�L�E��d�e�e�d�g��W��Y���W��^�D��d�e�w�u�w�}�B��D���V��^�D��e�d�y�`�`�`�W��I����V��_�E���`�m�h�u�f�l�F��H����V��NךU���l�u�k�w�g�l�F��H����W�X�U��w�e�d�d�g�m�F��I���W�	N��E��d�d�e�e�f�m�[�ԜY����F�L�D��e�d�e�d�f��W��Y���V��_�E��d�d�w�u�g�}�I���I����W��^�E���u�u�u�c�b�`�W��H����W��_�E���c�c�h�u�f�l�F��I����W��N�B��u�d�d�d�g�l�G��H���9F�X�U��w�e�d�e�g�l�G��H���_�	N��E��e�e�e�d�f�m�[��I���W��^�D��d�d�e�y�]�}�W��Y���V��_�D��e�e�w�u�f�}�I���I����V��^�E���u�d�u�k�u�m�F��H����V��B��U���c�a�h�u�f�l�G��I����V��N�@��u�d�d�e�g�m�F��H���W��
P��D��e�d�d�e�g�m�U���Y���Q�	N��E��e�d�e�d�f�l�[��A���W��^�E��d�d�d�y�a�d�J���H����V��^�D��y�_�u�u�e�}�I���I����W��^�E���u�g�u�k�u�m�F��I����V��B��G���k�w�e�d�g�m�G��H���l�N�F��u�d�d�d�f�m�F��I���T��
P��D��d�d�d�e�f�m�U���K���D��^�D��d�e�e�w�w�}�W��O���W��_�D��d�d�d�y�a�j�J���H����V��_�D��y�c�m�h�w�l�F��I����V��L����u�g�u�k�u�m�G��H����W��B��F���k�w�e�e�g�l�G��H���P��S�W��e�e�e�e�g�m�G��s���U��
P��D��d�d�e�e�f�l�U���J���D��^�E��d�e�d�w�w�n�W���[����V��_�E��w�u�u�u�a�h�J���H����V��^�D��y�c�c�h�w�l�F��H����W��L�C��h�u�d�d�g�l�G��H����FǻN��F���k�w�e�e�f�m�G��H���P��S�W��e�d�e�e�g�l�G��O���F�_�D��d�d�d�e�{�W�W���M���D��^�E��d�e�e�w�w�i�W���[����W��_�E��w�u�a�u�i��G��I����W��_��U���u�c�a�h�w�l�F��H����W��L�C���h�u�d�d�g�l�F��I����F��N��U��d�e�d�e�f�l�G���Y���P��S�W��e�e�d�e�f�m�G��O���F�_�E��e�e�e�d�{�k�N��Y����V��_�E��e�y�_�u�w�h�W���[����V��^�D��w�u�`�u�i��G��H����W��^��U���u�k�w�e�f�l�F��H����J�N��C��h�u�d�e�f�l�F��I����F��N��U��e�d�d�e�g�l�F���Y����X�^�D��d�e�d�d�u�}�W���O���F�^�D��e�e�d�e�{�k�@��Y����W��_�E��d�y�c�m�j�}�F��H����V��^�Y�ߊu�u�`�u�i��G��I����W��^��U��u�k�w�e�f�m�F��H����J�_��K���e�d�e�e�g�l�F��U���F��N��U��e�d�d�e�f�m�F���Y����X�^�D��d�d�d�e�u�}�A���G����W��_�D��e�w�u�u�w�k�B��Y����W��_�D��d�y�c�c�j�}�F��H����V��_�Y��b�h�u�d�g�m�F��I����D�=N��U��u�k�w�e�f�l�F��H����J�W��K���e�d�d�e�f�m�F��U����[�_�D��e�d�d�d�g�q�}���Y����X�^�E��e�e�e�d�u�}�@���G����W��_�E��d�w�u�b�w�c�U��H����V��^�W���u�u�c�a�j�}�F��I����W��^�Y��`�h�u�d�g�m�G��I����D�Y�H���d�e�e�d�f�m�F��[��ƹF� Y��K���e�d�e�d�f�l�G��U����[�_�D��d�e�e�d�f�q�A��D���V��_�E��d�e�y�_�w�}�O���G����W��^�D��d�w�u�m�w�c�U��H����W��_�W���m�u�k�w�g�l�G��H����W�d��U��f�h�u�d�g�m�G��I����D�V�H���d�e�e�e�f�l�G��[����F�L�E��e�e�d�d�f��W���Y����[�_�E��d�d�d�d�f�q�A��D���V��_�D��d�d�y�c�o�`�W��I����V��_�D���_�u�u�m�w�c�U��I����V��_�W���l�u�k�w�g�m�F��H����V�X�U��w�e�e�d�g�m�G��I���F�W�H���d�e�d�e�f�l�F��[���� F�L�E��e�e�e�e�g��W��Y���V��_�D��d�e�w�u�w�}�A��D���V��^�E��e�d�y�c�a�`�W��I����V��_�E���c�b�h�u�f�m�F��H����V��NךU���l�u�k�w�g�m�G��I����V�X�U��w�e�e�e�f�l�G��H���V�	N��E��e�e�d�d�g�l�[�ԜY����F�L�E��d�d�d�d�f��W��Y���V��^�E��d�d�w�u�g�}�I���I����V��^�E���u�u�u�b�c�`�W��I����W��_�E���b�`�h�u�f�m�F��I����W��N�C��u�d�e�d�g�m�F��H���9F�Y�U��w�e�e�e�g�l�F��H���^�	N��E��e�e�e�d�f�m�[��@���W��_�E��e�d�e�y�]�}�W��Y���V��^�E��e�e�w�u�f�}�I���I����W��^�E���u�d�u�k�u�m�G��H����V��B��U���b�f�h�u�f�m�G��I����V��N�A��u�d�e�e�f�l�F��H���W��
P��D��e�d�d�d�g�l�U���Y���P�	N��E��d�e�d�d�f�m�[��N���W��^�E��d�d�d�y�`�e�J���H����V��_�E��y�_�u�u�f�}�I���I����W��_�D���u�g�u�k�u�m�G��H����V��B��G���k�w�e�e�f�l�F��I���l�N�G��u�d�e�e�g�m�G��I���T��
P��D��e�e�d�e�f�m�U���K���D��^�E��d�e�d�w�w�}�W��L���W��^�E��e�d�e�y�`�k�J���H����V��_�E��y�b�b�h�w�l�G��I����V��L����u�g�u�k�u�m�G��H����W��B��G���k�w�e�e�g�l�G��H���Q��S�W��e�e�d�d�f�l�F��s���U��
P��D��e�d�e�e�f�m�U���J���D��^�D��e�d�e�w�w�n�W���[����V��_�E��w�u�u�u�`�i�J���H����W��^�D��y�b�`�h�w�l�G��H����W��L�B��h�u�d�e�g�l�G��I����FǻN��F���k�w�e�e�g�m�F��H���Q��S�W��e�e�e�e�g�m�G��N���F�^�E��e�e�d�d�{�W�W���M���D��^�E��d�e�d�w�w�i�W���[����V��_�E��w�u�a�u�i��G��I����V��^��U���u�b�f�h�w�l�G��I����V��L�B��h�u�d�e�g�m�G��I����F��N��U��e�e�e�e�g�m�F���Y���Q��S�W��e�e�d�e�g�m�G��N���F�^�E��e�d�e�e�{�j�O��Y����V��_�D��e�y�_�u�w�i�W���[����V��_�D��w�u�`�u�i��G��I����V��^��U���u�k�w�e�g�m�G��H����J�N��B��h�u�d�e�g�m�F��H����F��N��U��e�e�e�d�g�l�F���Y����X�^�E��e�d�d�e�u�}�W���N���F�^�E��d�e�e�e�{�j�A��Y����V��^�D��d�y�b�b�j�}�F��I����V��_�Y�ߊu�u�`�u�i��G��I����W��^��U���u�k�w�e�g�m�G��H����J�^��K���e�e�e�e�g�m�F��U���F��N��U��e�e�e�e�g�l�F���Y����X�^�E��e�e�e�d�u�}�A���G����V��^�E��d�w�u�u�w�j�C��Y����V��^�E��e�y�b�`�j�}�F��I����V��_�Y��c�h�u�d�g�m�G��I����D�=N��U��u�k�w�e�g�m�G��I����J�V��K���e�e�e�e�g�m�G��U����[�_�E��e�e�e�e�f�q�}���Y����X�^�E��e�e�e�d�u�}�@���G����V��^�E��d�w�u�b�w�c�U��I����V��^�W���u�u�b�f�j�}�F��I����V��_�Y��a�h�u�d�g�m�G��I����D� Y�H���d�e�e�e�g�m�F��[��ƹF� X��K���e�e�e�e�g�m�F��U����[�_�E��e�e�d�e�g�q�@��D���V��^�E��d�e�y�_�w�}�@���G����V��^�E��d�w�u�m�w�c�U��I����W��^�W���m�u�k�w�g�m�G��H����V�d��U��g�h�u�d�g�m�G��H����D� V�H���d�e�e�e�f�m�F��[����F�L�E��e�d�e�d�f��W���Y����[�_�E��e�e�d�e�g�q�@��D���V��^�D��e�e�y�b�`�`�W��I����W��_�E���_�u�u�m�w�c�U��I����W��_�W���m�u�k�w�g�m�G��I����V�Y�U��w�e�e�e�f�m�G��I���F� W�H���d�e�e�e�g�m�G��[����F�L�E��e�e�d�e�f��W��Y���V��^�D��e�e�w�u�w�}�@��D���V��^�E��e�e�y�b�b�`�W��I����W��^�D���b�c�h�u�f�m�G��H����W��NךU���l�u�k�w�g�m�G��I����W�Y�U��w�e�e�e�g�m�G��I���
_�	N��E��e�e�d�e�f�l�[�ԜY����F�L�E��d�e�d�e�f��W��Y���V��^�D��d�e�w�u�g�}�I���I����V��^�D���u�u�u�m�d�`�W��I����W��^�D���m�a�h�u�f�m�G��I����V��N�@��u�d�e�e�f�m�G��I���9F�V�U��w�e�e�e�f�l�F��H���Q�	N��E��e�d�e�e�f�m�[��A���W��^�D��d�d�e�y�]�}�W��Y���V��_�E��e�d�w�u�f�}�I���I����V��_�D���u�d�u�k�u�m�G��I����W��B��U���m�g�h�u�f�m�G��H����W��N�F��u�d�e�e�g�l�G��I���W��
P��D��e�e�e�e�g�m�U���Y���S�	N��E��d�d�d�e�g�l�[��O���W��^�D��e�e�d�y�o�j�J���H����V��_�D��y�_�u�u�f�}�I���I����W��_�D���u�d�u�k�u�m�G��I����W��B��G���k�w�e�e�f�m�F��H���l�N�D��u�d�e�e�f�l�F��H���T��
P��D��e�d�d�d�g�l�U���K���D��^�D��d�d�e�w�w�}�W��M���W��^�D��d�e�d�y�o�h�J���H����W��^�E��y�m�c�h�w�l�G��I����V��L����u�g�u�k�u�m�G��I����W��B��G���k�w�e�e�g�m�G��H���^��S�W��e�e�e�d�f�l�F��s���U��
P��D��d�e�e�d�g�l�U���J���D��^�E��d�e�d�w�w�n�W���[����V��^�D��w�u�u�u�o�n�J���H����W��^�D��y�m�a�h�w�l�G��H����W��L�M���h�u�d�e�f�l�F��H����FǻN��F���k�w�e�e�g�m�F��I���^��S�W��e�e�d�d�g�l�F��A���F�^�E��e�e�e�e�{�W�W���J���D��^�D��d�e�e�w�w�i�W���[����W��_�D��w�u�a�u�i��G��H����V��_��U���u�m�g�h�w�l�G��I����W��L�M��h�u�d�e�f�m�G��I����F��N��U��e�d�e�d�f�l�F���Y���^��S�W��e�d�e�e�g�l�G��A���F�^�D��d�e�e�e�{�e�@��Y����W��_�D��d�y�_�u�w�i�W���[����W��^�D��w�u�a�u�i��G��H����W��_��U���u�k�w�e�g�l�F��H����J�N��M��h�u�d�e�g�m�G��H����F��N��U��e�e�e�d�f�m�G���Y����X�^�E��e�e�e�e�u�}�W���A���F�^�E��d�e�e�d�{�e�B��Y����V��_�E��d�y�m�c�j�}�F��I����W��_�Y�ߊu�u�`�u�i��G��I����W��^��U���u�k�w�e�f�m�F��I����J�W��K���e�d�e�d�f�l�G��U���F��N��U��e�e�d�d�g�l�G���Y����X�^�E��e�e�d�e�u�}�A���G����W��^�D��e�w�u�u�w�e�D��Y����V��^�E��d�y�m�a�j�}�F��I����V��_�Y��`�h�u�d�g�m�F��I����D�=N��U��u�k�w�e�f�l�G��H����J�Y��K���e�d�d�e�f�m�F��U����[�_�D��d�d�d�e�f�q�}���Y����X�^�E��d�e�d�d�u�}�@���G����W��^�E��d�w�u�b�w�c�U��H����V��^�W���u�u�m�g�j�}�F��H����W��^�Y��f�h�u�d�g�l�G��H����D�Y�H���d�e�d�d�g�l�G��[��ƹF� [��K���e�d�e�e�g�l�F��U����[�_�D��d�e�d�d�f�q�O��D���V��_�E��d�e�y�_�w�}�@���G����W��^�E��e�w�u�b�w�c�U��H����V��_�W���m�u�k�w�g�l�F��I����V�d��U��d�h�u�d�g�l�G��I����D�V�H���d�e�d�d�g�m�F��[���� F�L�E��d�d�e�e�g��W���Y����[�_�D��d�e�d�d�g�q�O��D���V��_�E��e�e�y�m�a�`�W��H����V��_�E���_�u�u�m�w�c�U��I����V��^�W���m�u�k�w�g�m�G��I����W�V�U��w�e�e�e�f�m�F��I���F�W�H���d�d�e�d�g�l�F��[����F�L�D��d�d�e�e�f��W��Y���V��^�E��d�e�w�u�w�}�O��D���W��_�D��d�d�y�m�c�`�W��H����V��^�D���m�`�h�u�f�l�G��H����V��NךU���l�u�k�w�g�m�F��H����V�V�U��w�e�e�d�g�m�G��I���
^�	N��E��d�e�e�d�f�m�[�ԜY����
F�L�D��d�e�d�d�g��W��Y���V��_�D��d�e�w�u�g�}�I���I����V��^�D���u�u�u�l�e�`�W��H����W��^�E���l�f�h�u�f�l�F��I����W��N�A��u�d�d�d�f�m�G��H���9F�W�U��w�e�e�e�g�m�G��I���P�	N��E��e�d�e�d�f�m�[��N���W��_�D��e�d�d�y�]�}�W��Y���V��_�E��e�e�w�u�g�}�I���I����V��_�E���u�d�u�k�u�m�G��H����W��B��U���l�d�h�u�f�l�F��I����V��N�G��u�d�d�d�f�l�G��I���
W��
P��D��d�d�e�d�f�m�U���Y���R�	N��E��e�e�e�e�f�l�[��L���W��^�E��e�e�e�y�n�k�J���H����V��^�E��y�_�u�u�f�}�I���I����W��_�D���u�d�u�k�u�m�F��I����W��B��D���k�w�e�d�g�l�G��H���l�N�E��u�d�d�e�f�l�G��I���
T��
P��D��e�e�e�d�g�l�U���K���D��_�E��e�e�e�w�w�}�W��J���W��^�D��e�e�e�y�n�i�J���H����W��^�D��y�l�`�h�w�l�F��H����V��L����u�g�u�k�u�m�F��H����W��B��G���k�w�e�d�g�m�G��H���_��S�W��d�e�e�d�g�m�F��s���
T��
P��D��d�e�d�e�f�l�U���J���D��_�D��d�e�d�w�w�n�W���[����V��_�D��w�u�u�u�n�o�J���H����W��^�D��y�l�f�h�w�l�F��I����W��L�L��h�u�d�d�f�m�F��H����FǻN��F���k�w�e�d�f�l�G��H���_��S�W��d�d�e�e�f�m�G��@���F�_�D��d�d�d�d�{�W�W���J���D��_�D��e�d�e�w�w�n�W���[����V��^�D��w�u�a�u�i��F��I����V��_��U���u�l�d�h�w�l�G��I����W��L�L��h�u�d�e�g�l�G��H����F��N��U��e�e�d�d�f�l�G���Y���_��S�W��e�e�d�e�g�m�F��@���F�^�D��d�d�e�d�{�d�A��Y����V��^�E��d�y�_�u�w�i�W���[����W��_�E��w�u�a�u�i��F��H����W��_��U��u�k�w�d�g�l�F��I����J�N��L��h�u�d�e�g�l�F��H����F��N��U��e�d�e�d�g�m�G���Y����X�_�D��e�e�e�d�u�}�W���@���F�^�E��d�d�d�e�{�d�C��Y����W��_�D��e�y�l�`�j�}�F��H����W��^�Y�ߊu�u�`�u�i��F��H����V��_��U���u�k�w�d�g�l�G��H����J�V��K���d�e�d�d�g�l�G��U���F��N��U��e�d�d�e�g�l�F���Y����X�_�D��e�e�e�e�u�}�A���G����V��_�D��d�w�u�u�w�d�E��Y����V��^�D��d�y�l�f�j�}�F��I����W��^�Y��a�h�u�d�g�m�G��H����D�=N��U��u�k�w�d�f�m�G��I����J�X��K���d�d�e�d�f�m�F��U����[�_�D��e�e�e�d�g�q�}���Y����X�_�E��d�d�e�e�u�}�A���G����W��_�E��d�w�u�b�w�c�U��H����W��_�W���u�u�l�d�j�}�F��I����V��_�Y��g�h�u�d�g�m�F��I����D�Y�H���d�e�d�e�f�m�F��[��ƹF� Z��K���d�d�e�d�f�l�G��U����[�_�D��e�e�d�e�g�q�N��D���V��_�D��e�e�y�_�w�}�@���G����W��_�E��e�w�u�b�w�c�U��H����W��^�W���b�u�k�w�f�l�F��I����W�d��U��e�h�u�d�g�l�G��I����D�V�H���d�e�d�d�f�m�F��[����F�L�E��d�e�d�e�g��W���Y����[�_�E��e�e�e�e�f�q�N��D���W��^�D��d�e�y�l�b�`�W��H����W��_�D���_�u�u�m�w�c�U��I����W��_�W���m�u�k�w�f�m�G��I����V�W�U��w�d�e�e�f�l�F��I���F�V�H���d�d�e�e�f�l�F��[����F�L�D��e�e�d�d�g��W��Y���W��_�E��e�d�w�u�w�}�N��D���W��_�E��d�d�y�l�d�`�W��H����W��_�D���l�a�h�u�f�l�F��H����W��NךU���l�u�k�w�f�m�G��H����V�W�U��w�d�e�e�g�m�F��I���
Q�	N��D��e�e�d�e�f�m�[�ԜY����F�L�D��d�d�d�d�f��W��Y���W��_�E��e�e�w�u�g�m�J���H����V��_�E��y�_�u�u�g�l�J���H����V��_�D��y�d�e�u�i��F��H����V��^��U��f�h�u�d�f�l�F��I����D�=N��U��a�h�u�d�f�m�G��I����D�^�U��w�d�d�e�f�m�F��I���V��
P��D��e�e�d�d�g�m�U���Y���V��
P��D��e�d�d�d�f�m�U���I���F�_�E��d�d�d�e�{�l�G���G����W��^�D��e�w�u�u�w�l�F���G����W��_�E��e�w�u�e�f�`�W��H����W��_�D���d�d�u�k�u�l�F��I����W��B��U���d�d�u�k�u�l�F��H����W��B��E��h�u�d�d�f�m�G��I����F��[��K���d�d�e�e�f�m�F��U���F��X��K���d�d�e�d�g�l�G��U����F�L�D��d�d�e�e�g��W��A���W��_�D��e�e�e�y�]�}�W��@���W��_�E��d�e�d�y�f�o�W���[����W��_�D��w�u�e�d�j�}�F��H����W��^�Y�ߊu�u�e�g�j�}�F��H����W��_�Y��g�u�k�w�f�l�F��I����W�_�A��u�e�e�e�g�m�G��I���lǑV�����0�� ����(���0����l4��x8��U���!�<�2�_�2�4�W�Զ����J9��T��*���'�
�o�%�8�8��������l��P��U���u�4�1�e�#�-�K�������9K��N �����u�'�;�9�#���ԜY���Z �t!��*�����}�1�%�t�Iϳ�����VK�������u�u�u�u�w�9�߁����N��_��U��r�r�n�u�w�}����Y���F�N�����e�!�%�i�w�9���Y����������,�!�0�<�w�/��������9�������n�_�0�:�.�<����&����W9�������u�4�1�d�w�?����Y�����E_�����h�4�1�d�]�p��������G��D�����3�u�u�u�>�}�4���&����t#��V
��D���u�0�
�<�2�l�W������F�N�����d�!�%�i�w�2����Y���A�=N��U���9�0�_�u�w�}�W�������l��R�����d�_�u�u�w�3�W���s�˿�]��D�����&�4�0�:�]�3�W�������9l��E�����&�o�%�:�2�.�_���P����V��d��Uʼ�u�6�>�0�2�)�������A��N���ߊu�u�u�u�1�u����Y�����YNךU���u�u�u�u�g�a�W���Q����l/��r)��]���'�
�8�|�l�W�W���Y�Ʃ�WF��d��U���u�<�u�6�f�`�P���Y����l�N��U���u�$�u�h�:�0�4���&����t#��V
��D���%�|�u�u�w�}�Wϻ�ӏ��9F���U���_�;�u�'�4�.�L����ƾ�_]Ǒ="�����u���_�$�}�2���
����\��h_�AĴ�9�_�0�!�#�}�Gݚ�O�Ҋ�lV��h_�����
�u�&�u�w�:������ƹF�N�����<�!�u�u���2���D����9F�N��U���'�&��;�2�g�>���>���F��[�U���u�u��1�2�.����Y�ƅ�g#��eN�U��n�u�u�%�%�}�}���Y���A��CN�<����
���l�}�W���YӅ��\��yN��1�����_�u�w�}�W�������\��yN��1��������u����
����G�_��:����e�n�u�w�}�WϽ�I����}F��s1��2���_�u�u�u�w�m�Mϑ�-ӵ��l*��~-��0�����!��3�5�Z��=����|F��d��U���u�4�1�0�$�}�W���*����|!��h8��!����1�0�&�>�)�W���Y����g)�UךU���u�u�0�u�w��$���5����l�N��Uʤ�u�u� �u���8���&����|4��V�����u�u�u����G���s����V��C����=�!�6� �2�<����Ӌ��wV��(��E���d�
�4�'�f�4�}���Y����\��CN��G��f��
�
��l����&¹��^F��=N��U���u�:�!�}�w�}�W���Y����_�'��&������_�w�}�W���Y�ƭ�W��N��U���
���
��	�%�ԜY���F�N��E���u��
���L���Y���F��Oʚ�������!���6��ƹF�N��U���1�'�u�u���3���>����v%��eUךU���u�u�u�u�2�}�W���*����|!��d��U���u�u�u�$�w�}�"���-����t/��a+��:���_�u�u�;�w�2������Ɠ9l��P��U���8�g�e�f���(���H����A9��E�� ��u�:�%�;�9�}�Gݚ�O�Ҋ�lV��h_�����
�
�:�_�w�}�������9F�N��U���u�k�6�>�]�}�W���Y����F������e�_�u�u�w�}����GӅ��l�N��Uʤ�u�k�$�y�w�}�W�������[�V
�����y�u�u�u�w�>�F��Y����9F�N��U��h�u�d�n�]�3�W�������G��dװ