-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�g�e�f����(�����A�=N��U���6�>�o��w�	�(���0��ƹF��G1�����u��
���L���YӇ��@��CN�<����
���l�}�WϿ�&����\��b:��!�����n�u�w�<�(�������f2��c*��:���n�u�u�4��8����Y����`2��{!��6�ߊu�u�;���<����&����	F��=��*����
����u�FϺ�����O��N������'�;�0�n�8�F��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����E����o��u����>��Y����]9��{	�����
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���)����Z��1��D���u��
���(���-��� W��X����n�u�u�<��)����&ù��F��~ ��!�����
����_������\F��d��Uʼ�
�'�1�-�2�)��������	F��=��*����
����u�FϺ�����O��N������`�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�������/��d:��9�������w�n�W������]ǻN�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W�������G��h_��U���u��
����2���+������Y��E��u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�V�����;�f�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������z(��c*��:���u�n�0�1�]�W��������A��R��U���8�g�e�f���(���Kӏ��9F������!�4�
�:�$�����&����`2��{!��6��u�d�n�u�w�>�����ƭ�l��D�����
�u�u����>���D����l�N�����;�u�%���)�(���&����`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�E��w�_�u�u�8�.��������l��h��*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V�=N��U���&�4�!�4��	��������\��c*��:���
�����d��������\�^�E��e�e�e�e�g�m�G��Y����\��V ������&�`�3�:�i�Mύ�=����z%��r-��'���l�1�"�!�w�t�M���I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�����`�o�����4���:����W��S�����|�o�u�e�g�m�G��I����V��L�U���6�;�!�;�w�-�$���Ĺ��^9��N��1��������}�F�������V�S��E��e�e�e�e�g�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�e�e�w�]�}�W���
������d:��ӊ�&�
�u�u���8���&����|4�W�����:�e�u�h�u�m�G��I����V��^�W�ߊu�u�:�&�6�)����-����9��Z1�Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�l�G��I����l�N�����;�u�%���)�F�������	F��s1��2������u�f�}�������	[�^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�g�3�:�l�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��e�e�w�_�w�}��������C9��h��F���8�d�u�u���8���&����|4�W�����:�e�u�h�u�m�G��H����V��^�W�ߊu�u�:�&�6�)����-����9��Z1�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����]ǻN�����4�!�4�
��.�Fځ�
����\��c*��:���
�����d��������\�^�E��e�e�e�e�g�m�G��Y����\��V ������&�d�
�$��B��*����|!��h8��!���}�l�1�"�#�}�^��Y����W��^�E��e�e�e�n�w�}��������R��c1��D݊�&�
�c�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��^�E��u�u�6�;�#�3�W���*����^��D��B��������4���Y����W	��C��\��u�e�d�e�g�m�G��I����D��N�����!�;�u�%����������F��d:��9�������w�l�W������F��L�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�e�1�0�F���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�e�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�d�d�o���;���:����g)��^�����:�e�u�h�u��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������rF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EU��tN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��_�E��u�u�6�;�#�3�W�������l
��1��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�D��n�u�u�6�9�)����	����@��A]��D���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�e�e�e�e�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�F��I����V��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�
�#�g�`�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�l�F��Y����\��V �����:�&�
�#�e�l�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(ܘ�I����\��c*��:���
�����l��������\�^�D��d�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EU��+��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�D���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Nӂ��]��G��H���e�e�e�e�l�}�WϽ�����GF��h�����#�f�e�o���;���:����g)��\����!�u�|�o�w�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*��e�o�����4���:����W��S�����|�o�u�d�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���L����F��d:��9�������w�l�W������F��L�E��e�e�e�e�g�f�W�������R��V�����
�#�
��m��3���>����v%��eN��U���;�:�e�u�j��F��H���9F������!�4�
�:�$�����L���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����d�
�e�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��L�U���6�;�!�;�w�-��������9��N�&���������W��Y����G	�N�U��e�d�e�e�g�m�G��Y����\��V �����:�&�
�#�g�m�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����V��UךU���:�&�4�!�6�����&����lU��q(��U���
���
��	�%���Nӂ��]��G��H���d�d�d�d�f�l�F��H��ƹF��X �����4�
�:�&��+�O���Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��d�d�d�w�]�}�W���
������T�����d�
�u�u���8���&����|4�Y�����:�e�u�h�u�m�G��I����V��_�����u�:�&�4�#�<�(���
���� T��q-�E��o������!���6���F��@ ��U���o�u�e�d�f�l�F��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�d�w�]�}�W���
������T�����f�
�g�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�e�g�f�W�������R��V�����
�#�
�u�w�	�(���0����p2��F����!�u�|�o�w�m�F��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���a�1�"�!�w�t�M���I����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�a�3�*����P���V��^�����u�:�&�4�#�<�(���
����9��N��1��������}�CϺ�����O�
N��E��w�_�u�u�$�:����	����U��N��1��������}�F�������V�S��E��e�e�e�e�g�m�G��[���F��C�� ���3�8�0�6�3�3�W�������l�N����� �0�3�8�2�>����Y����C9��h��U���<�;�9�<�w�3����s���@��V�����2�6�0�
��.�F������5��h"��<��u�u�&�2�6�}��������lU��N��:����_�u�u�>�3�Ͻ�&����q'��X�� ���b�e�0�e�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�L���Yӕ��]��T��0����� �%�#�n�(߁�&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����4�u�'�
�"�l�F���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����d�b�o����0���/����aF�N�����u�|�_�u�w�4��������T9��R��!���f�3�8�g�m��3���>����F�D�����%�&�2�7�3�k�W���6����}]ǻN�����9�4�
�<��.����&����U��N�&������_�w�}����Ӈ��@��U
��B���u����l�}�Wϭ�����T��Q��F݊�g�o�����4���:����U��S�����|�_�u�u�>�3�Ϭ�����\��c*��:���
�����l��������l�N�����u�%�&�2�4�8�(���
�ғ�@��T��!�����n�u�w�.����Y����Z��S
��M������]�}�W�������V�� V��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�'�.��������l��1����o������}���Y����R
��G1�����1�l�u�u���6��Y����Z��[N��*���
�&�$���)�A�������	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������@��1�����0�1�3�
�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��[1��0����:�!� ��j����H����_��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��%�"�������R��h��F���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����2��x��Mފ�
�0�
�g�`�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h]�����e�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y���� R��R	��G��o������!���6�����Y��E��u�u�&�2�6�}�$���,����|��[��*���`�e�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l��{:��:���c�
�
�0��o�@��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����&�����!�d�o�;�(��&���5��h"��<������}�f�9� ���Y����F�D����������)�F�������Q��N��1��������}�D�������V�=N��U���;�9�4�
�>�����*����9��Z1�Oʆ�����]�}�W�������C9��P1����l�o�����}���Y����R
��G1�����0�
��&�f�����I����g"��x)��N���u�&�2�4�w�-��������_�,��9���n�u�u�&�0�<�W���&�Г�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Cف�����
S�=��*����
����u�W������]ǻN�����9�!�%�`��(�O���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�g�'�2�f�m�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
�
� �m�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
�
�0�
�d�k�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����<�3�
�a��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����<�'�2�d�f�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Gӊ�
� �m�d�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Gӊ�
�0�
�f�o�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��B���3�
�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��B���'�2�d�g�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������_9��y*�����
�m�0�g�1��Bہ�J����g"��x)��*�����}�d�3�*����P���F��P ��U������!�%��O���K����lW��N�&���������W��Y����G	�UךU���<�;�9�4��4�(�������@��h��*��o������}���Y����R
��G1�����1�d�f�o���2���s���@��V��&��� ���!��1����&�ߓ�V��]�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�����
����g9��]�����g�o�����4�ԜY�ƿ�T�������7�1�d�g�m��8���7���F��P ��U�������#�h�(���@�Г� F��d:��9�������w�n�W������]ǻN�����9�4�
�<��.����&����l ��h_�Oʆ�����]�}�W�������C9��P1����g�o�����}���Y����R
��X������!�a�
�"�l�F߁�K����g"��x)��*�����}�u�8�3���B�����Y�����
��,� ��e����H����	F��s1��2������u�g�9� ���Y����F�D�����%�&�2�6�2��#���HĹ��^9��T��!�����n�u�w�.����Y����Z��S
��E���u����l�}�Wϭ�����U5��r"��!���
�e�
�
�"�d�O���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�
�f�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��D���%�u�u����>���<����N��
�����e�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�4�
�<��.����&����l ��h_�Oʆ�����]�}�W�������C9��P1����g�o�����}���Y����R
��E�� ��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U��Y��D��������4���Y����W	��C��\�ߊu�u�<�;�;�:����&����CV�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�l�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����a�
� �d�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��Aފ� �d�l�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����G��Y�� ��a�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��B1�A���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������
9��T��!�����
����_������\F��d��Uʦ�2�4�u�9���5�������G9��h��*ۊ� �d�d�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������`9��u;��9���'�
�g�3��m�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
� �g�g�-�W���-����t/��a+��:���b�1�"�!�w�t�}���Y����R
��X��*ي� �g�e�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����G��^1����
� �g�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��*��� �g�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V��h��*���g�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��1�����3�
�a�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���3�
�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���3�
�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����A��1�����6�&�
�4�#�;�(��&���5��h"��<������}�c�9� ���Y����F�D�����0�
�8�
�e�;�(��&���5��h"��<������}�c�9� ���Y����F�D�����
�0� �!�a����O����	F��s1��2������u�f�}�������9F������3�
���e����&����K��h_�� ��a�%�u�u���8���&����|4�Y�����:�e�n�u�w�.����Y����Z9��h]�*��o������!���6�����Y��E��u�u�&�2�6�}����Iƹ��U��X��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�d����O����	F��s1��2������u�`�9� ���Y����F�D�����8�
�`�3��n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �f�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������\��D���3�
�d�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hY�����
�a�
�f�m��3���>����v%��eN��Eʱ�"�!�u�|�]�}�W�������l4��B��Cۊ� �f�a�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��z;��G���!�m�
�;�1�	��������l��N��1��������}�F�������V�=N��U���;�9�&�9�#�-�(�������l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�j����&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'��(���J�ԓ�F��d:��9�������w�m��������l�N�����u��-� ��3����M���� P��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�8�1����&����CT�=��*����
����u�W������]ǻN�����9�%��9�����A����	F��s1��2������u�d�}�������9F������9�6��3��l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����d�3�
�g��l�Mύ�=����z%��r-��'���g�1�"�!�w�t�}���Y����R
��Z��*���a�3�
�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�����
�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƾ�G9��Q��FҊ�f�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	����l��h��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��Q��CҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l��B1�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����H����R��T��*���a�g�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�_9��G1�����c�
�f�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��V��C1�����m�
�f�o���;���:����g)��_����!�u�|�_�w�}����Ӏ��K+��c\�� ���`�<�
�-���(���M�Г�F��d:��9�������w�l�W������]ǻN�����9�!�%�&�1��G݁�K����g"��x)��*�����}�u�8�3���B�����Y�����g�
� �`�o�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��M���
�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��@���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��X��D��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�%�e�g��(���L�֓� F��d:��9�������w�o�W������]ǻN�����9�!�%�g��(�B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ��&�9�
�n�;�(��&���5��h"��<������}�f�9� ���Y����F�D������-� ��9�(�(�������g��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������C9��h[�*��o������!���6�����Y��E��u�u�&�2�6�}�����ד�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����R��N�&���������W������\F��d��Uʦ�2�4�u��/��#ݰ�����l ��X�����u��
����2���+������Y��E��u�u�&�2�6�}�$���5����F��V�� ��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4����	����9��h��C���%�u�u����>���<����N��
�����e�n�u�u�$�:��������9��hX�*��o������!���6�����Y��E��u�u�&�2�6�}����&ƹ��lP��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-����&����lP��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��(�������U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%��1�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�:���(���O�ߓ�F��d:��9�������w�j��������l�N�����u�:�
�
��(�A���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʡ�%�<�<�
��(�A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
�d�<�1��Aց�K����g"��x)��*�����}�u�8�3���B�����Y�����9�
�g�3��e�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
� �c�b�-�W���-����t/��a+��:���b�1�"�!�w�t�}���Y����R
��X��*ӊ� �c�`�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����G��^1��*���c�3�
�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1��؊�
� �b�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������E��*���b�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӈ��_��h��B���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����l �� Z�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�3����K����U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�n�(���N�ߓ�F��d:��9�������w�m��������l�N�����u�8�
�m�1��C؁�K����g"��x)��*�����}�u�8�3���B�����Y�����f�
� �b�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E�� ��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������@U��B1�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�����Փ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�C݁�����l��N��1��������}�GϺ�����O��N�����4�u�8�
�d�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�a�
� �f�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��_�� ��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������_��R�����<�3�
�b��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�D���8�'�4�
��(�@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
� �m�f�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_�*���:�2�;�<�1��Dց�K����g"��x)��*�����}�u�8�3���B�����Y�����a�
� �b�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
�
�0�:�0�3����Kƹ��\��c*��:���
�����}�������9F������!�%�a�
�"�j�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�
�
�"�e�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�
�
�"�e�@���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�
�
�8����@����	F��s1��2������u�g�9� ���Y����F�D�����8�
�m�3��m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�m�<�3��h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �m�f�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[�����m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����v*��c!��*��
� �m�m�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��^��*��� �l�a�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����@��C��G���3�
�d�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��Gۊ�
� �l�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��[1�����<�3�
�g��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1�����d�g�g�3��d�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&���'�d�d�g�f�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����0�
�8�a�����M����	F��s1��2������u�d�}�������9F������&�9�!�%�g�4����M¹��\��c*��:���
�����l��������l�N�����u�0�
�8�b��(���@�ޓ� F��d:��9�������w�n�W������]ǻN�����9�3�
���	����A����
P��G^��U���
���
��	�%���Y����G	�UךU���<�;�9�3���3�������G	��Y�� ��a�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����P��B1�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����@¹��l_��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�9�)��������9��T��!�����
����_�������V�=N��U���;�9�;�!�?�i����@����\��c*��:���
�����}�������9F������!�%�`�
�"�l�Gہ�K����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$����������
F��d:��9����_�u�u�>�3�Ͽ�&����Q��Y�Oʗ����_�w�}����Ӗ��R
�� Z�� ��d�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӊ��l0��1��*��l�%�u�u���8���&����|4� N�����u�|�_�u�w�4��������lW��Q��E���%�u�u����>���<����N��
�����e�n�u�u�$�:��������ZW�� 1��*��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϭ�����U��Z�����u��
����2���+������Y��E��u�u�&�2�6�}����J¹��ZW��B1�@ي�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������ZT��T��*���!�3�
�e�n�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��D�����<�
� �d�a��D��*����|!��h8��!���}�a�1�"�#�}�^�ԜY�ƿ�T�������!�c�
� �f�d�(��Cӵ��l*��~-��0����}�b�1� �)�W���s���@��V��&��� ��;� ��o��������9��h_�F���u�u��
���(���-���Q��X����n�u�u�&�0�<�W���&�ӓ�F9��W��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������S��N�&���������W������\F��d��Uʦ�2�4�u�8��n����H�ד�F��d:��9�������w�m��������l�N�����u�8�
�a�1��F���	����`2��{!��6�����u�b�3�*����P���F��P ��U���
�e�3�
�f�n����Y����)��t1��6���u�b�1�"�#�}�^�ԜY�ƿ�T����*���3�
�d�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������_��D���
�d�b�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����G��Y�� ��`�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��V��C1�*���d�c�
�`�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��b"�����
�g�<�
�'�$����&����l��N��1��������}�F�������V�=N��U���;�9�&�9�#�-�(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'����Aƹ��\��c*��:���
�����}�������9F������&�9�!�%��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʳ�
���g��)�A݁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u����4�������9��h_�A���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���������C1�*؊� �d�l�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��D���6�u�u����>��Y����Z��[N��*���
�&�$���)�N�������	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������F9��1�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Mǹ��lW��h�����o������!���6�����Y��E��u�u�&�2�6�}����N����S��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����_��G����������4���Y����\��XN�N���u�&�2�4�w�-��������C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�<�;�;�<�(�������l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�&�2�6�}��������9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1��������lU��E��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�&�0�<�W���7����^F��d:��9�������w�l�W������]ǑN�����:�0�!�8�e�m�Dۘ�&ù��W�� ��Fػ�
�g�f�3�;�����*�����R��U�ߊu�u�u�u��g�>���>����F�N��;������o��	�0���s���F�S��*����u�u����L���Y�����1��1���o�����W�W���Y�ƨ�F��~*��U������u�l�}�WϮ����F�N�����o��u����>��Y���F��R��U���������}���Y���W��T��;ʆ�������8���J�ƨ�D��^����u�u�u�<�f�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Y�����N��U���
���n�w�}�W�������	F��cN��1��������}�D�������V�UךU���;�u�:�%�9�3�L�ԶY����\��Y��U���c�a�3�g�;����K������\��*���
�&�u��w�}�������9F�N��U���o�����W�W���Y�Ƃ�~9��v)��Oʜ����_�w�}�W����֓�z"��T��;����n�u�u�w�}����&����{F��~ ��2���_�u�u�u�w�2����=���/��r)��U��u�u�%�'�w�W�W���Y�ƨ�]V�'��&���������W��Y����G	�UךU���u�u�<�d�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����\��N��!ʆ�������8���J�ƨ�D��^��\�ߊu�u�;�u�8�-����B��ƹF��X�����u�e��c�c�;�G�������]�� ��D���_�u�u�2�8����s���F�~*��U�����n�u�w�}�Wϐ�4����t#�'��0���n�u�u�u�w�9�߁�0����	F��c+��'�ߊu�u�u�u�>�l� ���1����}2��r<�U���u�u�1� ���#���Y����t#��UךU���:�!�}�u�w�}�WϺ�����z(��c*��:���
�����l��������l�N��Uʱ�;�u�u����;���:����g)��]����!�u�|�_�w�}�W���	����\��yN��1��������}�CϺ�����O��N��U���1� �u�u��}�#���6����e#��x<��Eʱ�"�!�u�|�~�W�W����Ư�^��R ���ߠ7�2�;�u�w�;�G�������]�� ��F؊�
� �9�1�'��W�������V��Z^��E���
�
�4�3�n����K����9��Q��*���_�u�u�0�2�4�W���Y���F�N��U��d�_�u�u�w�}�"���-����X�d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�o�}���Y���W	��h9��!���k�f�|�u�w�-�������F�N�����h�u�%�6�<�W�W���Y�ƾ�@��
P�����!�_�u�u�w�}���D�ƫ�C9��h_�*��_�u�u�u�w�4�F��Y����U��_��D�ߊu�u�u�u�2�`�W���&���� W��RBךU���u�u�:�!�j�}��������l��dךU���
�
�8�9�d�3�(���
����9��O1�����u�u�:�%�9�3�W��=����u ��h����;�
�g�&�d��(���&����F�P�����8�%�}�u�w�}�Wϗ�Y���l�N��Uʛ�����j�}�[���Y�����1��1���h�u�g�_�w�}�W����ד�z"��S�F���u�u�u�u�3�(�(���-���U��=N��U���!�8�%�}�w�}�W�������X��E�� ��b�%�y�u�w�}�WϺ������h��D���%�y�u�u�w�}����Y����A��B1�B���|�_�u�u�1�m����&�Ԣ�lU��D1��D���u�u�:�%�9�3�W��=����u ��h����;�
�g�&�f�l�W�������Z��V�����u�u�u��j�}�[���Y���(��h=��2���k�d�_�u�w�}�W���I����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���:�!����`�W���Y����\��Z��]���u�u�u�1�9�}�IϹ�	����R��G^�U���u�u�1�;�w�c�������� 9��d��U���u�:�6�1�w�c�������� 9��T��Y���u�u�u�1�"�}�IϹ�	����R��G\����u�3�e�3�:��E���J����9��bY��U���%�;�;�u�g��A����֓�P��\��*���&�d�d�u�w�:����Ӌ��NǻN��U����h�u�y�w�}�W���7����g'��S�D�ߊu�u�u�u�>�m� ���1��� T�N��U���1�;�
���}�I��U���F�
�������h�u�~�}�WϮ��ơ�CF�N��U���1�;�u�k�#�-�Cہ�����l��=N��U���u�<�d�h�w�0�(�������
9��d��U���u�:�6�1�w�c����Mǹ��lW��h�����_�u�u�u�w�2���Y����R��B1�L���|�_�u�u�1�m����&�Ԣ�lU��D1��D���u�u�:�%�9�3�W��=����u ��h����;�
�g�&�f�l�W�������Z��V�����u�u�u��j�}�[���Y���(��h=��2���k�d�_�u�w�}�W���I����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���:�!����`�W���Y����\��Z��]���u�u�u�1�9�}�IϪ�	����U��Z��E�ߊu�u�u�u�>�l�J�������l ��[�����u�u�u�u�8�>����GӒ��lR��Q��@ފ�%�:�0�_�w�}�W������F��G1�*���d�a�%�|�]�}�Wϸ�I����C9��Y��G���d�d� �u�w�2�����ơ�"��Z��*ڊ�6�%�f�;��o����H�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�f�W�W���Y�ƨ�]V��~*��U��f�y�u�u�w�}����&����{F�]����u�u�u�:�#�
�3���D����9F���ʸ�%�}�u�u�w�}����Y����^��1��*���
�e�_�u�w�}�W���H���G��_�� ��l�%�y�u�w�}�Wϱ�����X��Z��D���
�`�
�%�8�8�}���Y���W	��S����`�
� �d�n�-�^�Զs��ƹF�N��ʶ�'�0�!�&�6�8�_���:����^O��QN��ʦ�4�0�8�6�>�8�W��Y����C9��h��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�%������DӇ��`2��C_�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�4��8����I����TF��D��U���6�&�{�x�]�}�W�������]9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�%�%�)����&����Z�V�����
�#�g�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���Kù��^9��G�����u�u�u�u�w�}�W���Y�����E�����
�'�2�i�w��$���:����lS��1��*��a�%�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��*��� �;�d�%�2�}����Ӗ��P��N����u�%�'�!�%��(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F������'�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��N���Y����l�N��U���u�u�u�u�w�<�(�������l��PN�U���
�b�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��*��� �;�g�%�2�}����Ӗ��P��N����u�%�'�!�%��(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F������'�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��N���Y����l�N��U���u�u�u�u�w�<�(�������l��PN�U���
�c�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��*��� �;�f�%�2�}����Ӗ��P��N����u�%�'�!�%��(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F������'�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��N���Y����l�N��U���u�u�u�u�w�<�(�������l��PN�U���-� ��;�"��E�������
Q��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�b�3�8�f�t�^Ϫ����F�N��U���u�7�:�
��$����A����lW�� N�U���9�-���#�i�(���H����CT��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�g�1�0�F���PӒ��]l�N��U���u�u�u�6���3�������9��1����f�u�h�6���3�������9��1��*���
�f�_�u�w�}�W���Y���P
��r+��4��� �%�!�f���(���DӀ��`#��t:����c�g�3�
�e��D�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h_��U���6�|�4�1�9�)�_���
����[��G1�����9�2�6�e�~�t����s���F�N��U���6�
������������9��N�U����
�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G��U���;�u�u�u�w�}�W���YӀ��`#��t:����m�'�2�d�`�}�Jϸ�&����p2��C1�M���
�e�
�f�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GR��D��\ʴ�1�;�!�}�9�/����M����W9��V
�� ��
�g�h�4��2����¹��O�C�����u�u�u�u�w�}�W���������C1�*؊�0�
�g�b�k�}�$���,����|��[��*���`�e�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� 9��Z1�\���=�;�u�u�w�}�W���Y����`9��b"�����
�a�d�'�0�l�B���DӀ��K+��c\�� ���a�d�3�
�o��D�ԜY���F�N��Uʡ�%�f�
�0��o�E��Y���� R��B1�G���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���J����lW��G�����u�u�u�u�w�}�W�������f*��x��8���<�9�
�l�%�:�F��Y����A��B1�B���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���J����lT���]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�}����Y���F�N��U���0�
�c�u�j�:����&����CT��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�b�1�0�A������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GR��D��\���u�=�;�u�w�}�W���Y�����h_�U��2�%�3�
�d��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Dڊ�&�
�|�u�%�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O�N���ߊu�u�u�u�w�}�W�������F�	��*���d�d�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����W��D��E���u�=�;�u�w�}�W���Y�����h��Dۊ�
�0�
�f�a�a�W���&����9��Q��Dӊ�g�_�u�u�w�}�W���Y�ƿ�_9��G\�����2�d�d�u�j�.����	�֓�l ��Z����u�u�u�u�w�}�W���
����^��h�����f�m�i�u�2����&����l^��h����u�u�u�u�w�}�W���&����9��E��D��u�h�&�9�#�-�@�������9��d��U���u�u�u�u�w�)���&����T��R�����a�
� �b�b�-�L���Y���F�N��U���
�g�'�2�f�m�W������9��hV�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����;�-�u�!�#�}����*����F����U���!�u�4�=�9�s�Z�ԜY�ƭ�l(��Q�����2�
�'�6�m�-����
�έ�l��E�����3�8�u�'�>�^���Yӄ��ZǻN��U���4�0�4�
��;�Ϸ�s���F�N�����u�%��
�#�����Y���F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u��������F��h�����:�<�
�|�~�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��D���8�e�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����9��Z1�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���g�3�8�d�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��[��U���u�u�u�u�w�}�W�������l ��R������&�f�3�:�o�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��A���8�f�h�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�c�;���s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���`�3�8�a�j�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!��.�(��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�B�������F�N��U���u�u�0�1�>�f�W���Y���F��_������&�c�3�:�h�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���O����lS��N��U���u�u�u�u�2�9���Y���F�N�����4�
��&�`�;���D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����l ��hX�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�O������FǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���@����l^�	NךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�4�
��1�0�K���	����@��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��L���8�m�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����V��D��U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��Dۊ�&�
�e�_�w�}�W���Y���F��DךU���u�u�u�u�w�}�W���	����U��S�����
�!�e�3�:�d�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��Dۊ�&�
�e�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�g�1�0�F��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Fށ�
����l�N��U���u�u�u�0�3�4�L���Y���F���ʴ�
��&�d��.�(��D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���J����lW��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��D��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���H����^9��S����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�4�
��;���Y����g9��Z�����f�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���f�3�8�d�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӈ��`2��C_�����d�u�k�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�d�
�&��i�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�i����H��ƹF�N��U���u�u�;�u�1�W�W���Y���F��R �����
�!�`�3�:�l�W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Fف�
����l�N��U���u�u�u�0�$�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����l ��h_����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��D��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��D܊�&�
�`�_�w�}�W���Y���F��SN��N���u�u�u�u�w�*����	����@��h��*��h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���m�3�8�d�l�}�W���Y���F������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�d��.�(��s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���d�
�&�
�`�`�W���Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�d����H��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���H˹��^9��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���;�4�
��$�l�(���&���FǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����l ��h_����u�u�u�u�w�}�W������F�N��U���u�u�u�%������DӇ��`2��C_�����d�n�u�u�w�}�W���Y����]��QUךU���u�u�u�u�?�3����-����9��Z1�U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��D���8�e�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�e�3�8�f�f�W���Y���F�N�����3�_�u�u�w�}�W�������G��DN��U�ߊu�u�u�u�w�}�W���	����U��S��-���������/���[���F�N��ʶ�&�n�u�u�2�9��������9F�C����:�0�4�&�0�}����
���l�N��*���0�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��*���u�%�&�2�4�8�(���
����U��W��U���7�2�;�u�w�}�WϷ�Y����\�V�����
�:�<�
�w�}���������F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�u�%�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������
O�N�����u�u�u�u�w�}�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�1�;�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�4����
������T��[���_�u�u�%�>�1�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�_�u�w�8��ԜY���F��F�����4�
�:�&��2����Y�ƭ�l��E��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������9F�N��U���u�%�<�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����0�1�u�&�>�3�������KǻN�����4�,�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����֓�@��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӇ��A��NN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����F��N�����u�'�6�&�y�p�}���Y����V��Y1�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�m����H����`9��{+��:���`�
�
� �f�m�(��Y����V��Y1�����|�u�u�7�0�3�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�l�|�u�?�3�}���Y���F�V�����;�e�i�u���;���6����9��Q��G���%�n�u�u�w�}����Y���F�N��U���'�!�'�
�w�`��������lV��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�/����&�ƭ�@�������{�x�_�u�w�-��������R��P �����o�%�:�0�$�<�(���Y����Q�������6�0�
��$�o�(���&���R��R�����%�0�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�l�~�}����s���F�N�����0� �;�d�k�}����N��ƹF�N�����_�u�u�u�w�}�W�������]9��S�����!�'�
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h�� ���g�4�&�2�w�/����W���F�V�����;�g�4�&�0�����CӖ��P����*��y�4�
�0�w�-��������`2��C\�����d�y�4�
�2�(����	����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����_�N�����u�u�u�u�w�}��������lT�
N����b�_�u�u�w�}����s���F�N�����0� �;�g�k�}��������9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��8����JӇ��Z��G�����u�x�u�u�6������Փ�@��Y1�����u�'�6�&��-�������T9��R��!���g�
�&�
�n�}�$���,����|��\��*���d�l�
�f�w�-��������C��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���=�;�_�u�w�}�W���Y����V��Y1�I����-� ��9�(�(���K����W��h����u�u�u�9�2�W�W���Y���F��h�� ���f�i�u�%�%�)����&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��G���
������T��[���_�u�u�%�$�:����H�Г�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��X��H���%�6�;�!�;�l�F������l ��_����!�u�`�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�a�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��Eʱ�"�!�u�e�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����N�ƭ�@�������{�x�_�u�w�-��������U��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��B���h�}�%�6�9�)����H����C9��h��]��1�"�!�u�f�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����g�1�"�!�w�o�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��\�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����l�u�h�}�'�>�����ד�[��G1��*���}�f�1�"�#�}�D���s���V��G�����_�_�u�u�z�<�(���&����V��V�����'�6�&�{�z�W�W���	����l��h\�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�e�u�h��-��������lW���6���&�}�c�1� �)�W��P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Gފ�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�g�u�j�u��������EW��S�����
�&�}�u�8�3���P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��F؊�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�f�u�j�u��������EW��S�����
�&�}�b�3�*����N����F�R �����0�&�_�_�w�}�ZϿ�&����Q��V�����;�%�:�0�$�}�Z���YӇ��@��U
��FҊ�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�i�w�<�(��������Y��E���u�%�6�;�#�1�F��B����������n�_�u�u�z�}��������lP�������%�:�0�&�w�p�W�������T9��S1�A���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�c�a�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��N�����u�'�6�&�y�p�}���Y����Z��S
��M���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�c�u�h��-��������lW���6���&�}�u�:�9�2�E���s���V��G�����_�_�u�u�z�<�(���&����Q��D��ʥ�:�0�&�u�z�}�WϿ�&����Q�� Y�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����b�i�u�4��2����¹��F��h-�����c�1�"�!�w�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����d�i�u�4��2����¹��F��h-�����d�u�:�;�8�l�^��Y����]��E����_�u�u�x�w�-��������F��D��U���6�&�{�x�]�}�W���
����W��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����u�h�}�%�4�3����H�����t=�����u�:�;�:�d�t�}���Y����C��R���ߊu�u�x�4��4�(���&����@��YN�����&�u�x�u�w�<�(���&����
^��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��M��u�4�
�:�$��ށ�Y�ƭ�l%��Q��Lʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����9��Z1����2�u�'�6�$�s�Z�ԜY�ƭ�l��h�����
�!�e�3�:�d��������\������}�%�&�2�5�9�N���Y����V��=N��U���u�3�}�%�$�:����@����[��=N��U���u�u�u�%�$�:����&����GW��Q��L��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��Dڊ�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����9��Z1�U���<�;�%�:�2�.�W��Y����C9��P1������&�d�
�$��G���
����C��T�����&�}�%�&�0�?���@���F��P��U���u�u�<�u�6���������
O��_�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�d�3�8�f�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C_�����d�u�&�<�9�-����
���9F������6�0�
��$�l�(���&�ד�@��Y1�����u�'�6�&��-��������U�N�����;�u�u�u�w�4�Wǿ�&����Q��Y�U���;�_�u�u�w�}�W���	����l��F1��*���g�3�8�d�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!�e�;���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���f�3�8�d�w�.����	����@�CךU���%�&�2�6�2��#���H����^9��h�����%�:�u�u�%�>����	����l��h_�\���u�7�2�;�w�}�W�������C9��P1����g�u�=�;�]�}�W���Y���R��^	������
�!�f�1�0�F���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$����������F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�a�1�0�F���
������T��[���_�u�u�%�$�:����&����GW��Q��Dي�&�<�;�%�8�}�W�������R��^	�����l�|�u�u�5�:����Y����������7�1�d�g�w�5��ԜY���F�N��*���
�&�$���)�C�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����l ��h_�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�A�������R��P �����&�{�x�_�w�}��������B9��h��C���8�d�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�e�~�}�Wϼ���ƹF�N�����%�&�2�7�3�l�A������F�N��U���4�
�<�
�$�,�$����Г�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��X�����`�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����ѓ�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�b�3�8�f���������PF��G�����4�
�<�
�3��G���Y����V��=N��U���u�3�}�%�$�:����K���G��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�c�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*��4�&�2�u�%�>���T���F��h��*���$��
�!�o�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lT��N�����u�u�u�u�w�}��������V��c1��DҊ�&�
�b�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�d�
�$��@��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��Dӊ�&�
�m�4�$�:�W�������K��N�����<�
�&�$����������9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��@���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��e�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�d�3�8�g�<����Y����V��C�U���4�
�<�
�$�,�$���¹��^9��V�����'�6�o�%�8�8�ǿ�&����Q��V��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��F���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�3�8�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�f�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�l�6�.��������@H�d��Uʴ�
�<�
�&�&��(���I����lW��V�����'�6�o�%�8�8�ǿ�&����Q��Y����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�g�
�$��N��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�E߁�
����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�f�3�:�o�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�\���u�7�2�;�w�}�W�������C9��P1����|�!�0�u�w�}�W���Y����C9��P1������&�f�3�:�o�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�n����K���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���a�3�8�f�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&���� 9��D��*���6�o�%�:�2�.��������W9��d��Uʷ�2�;�u�u�w�}��������T9��S1�\ʡ�0�u�u�u�w�}�W�������T9��R��!���a�3�8�f�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�a�1�0�D��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��@���8�a�4�&�0�}����
���l�N��*���
�&�$���)�(���&ǹ��@��h����%�:�0�&�6���������
OǻN�����_�u�u�u�w�;�_���
����W��W�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�a�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�`�3�:�i�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�����c�4�&�2�w�/����W���F�V�����&�$��
�#�����&����T��E��Oʥ�:�0�&�4��4�(���&���F�U�����u�u�u�<�w�<�(���&����Q�C��U���u�u�u�u�w�<�(���&����l5��D�����c�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���b�3�8�c�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��Q��Bʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�
�$��(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��1����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�b�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���7�:�
��.�(�(�������V��N�U¡�%�`�
� �f�m�(������A��B1�F���|�_�u�u�;��9�������^��h\�� ��a�%�u�h�]�}�W���Y����*��Y	��L���d�"�0�u�$�1����N����V��\�E���u�d�|�0�$�}�W���Y����V
��Z�*��� �l�m�%�l�}�WϽ�&����q'��X�� ���b�0�d�d�1��Nށ�I���V�^ �����
�y�:�=�%�`�P���B�����q+��7���:�!� �
�`�8�F�������9��R�����u�u�u�%�4�3����J����D��F��*������ �'�)�D؁�&¹��U��_��E��u�u�d�|�2�.�W���Y�����q+��7���:�!� �
�`�m���s���U5��r"��!���
�e�
�
�"�d�O���Y���F�N�������� ��i�(���&������YN�����8�f�
�
�2��D��I���W����ߊu�u�u�u�2����&����l_��h����u��������O����Q��G]��H�ߊu�u�u�u�'�>��������F��R �����f�
� �m�d�-�_���D����F��D��U���u�u�'�2�f�j�}���Y����v*��c!��*��
� �c�g�'�}�J���D͏��A��C1�U���0�&�k�x�~�W�W���*����v%��B��AҊ� �c�g�%�w�`�}���Y���U5��z;��G���!�c�
�
�2��E������ ��d+��6���!�d�m�3��m�(��I���W����ߊu�u�u�u�;��2���:����C��Y��*���n�u�u�3���2�������lT��B1�Eފ�f�i�u�u�w�}�WϹ�	����U��G\�����}�:�9�-�����&����U��^��H��r�u�9�0�]�}�W���Y����Q��=N��U�������#�h�(���@�Г�F�F�K���'�&�!�a�w�)����G���l�N��*����� �
�o�;�(��&���FǻN��U���%�6�;�!�;�n�(������U5��r"��!���
�m�3�
�a��G��Y���O��[�����u�u�u�;��<����I����l�N��*��� ���0�:�o�(���K�Г�F���%���4�;�
�
��f�W�������A��^��D���
�l�
�f�k�}�W���Y����]9��{�����
�
�u�=�9�u����I����^��G\��\��r�r�u�9�2�W�W���Y�ƾ�T9��UךU����!�'�d�f�o�E���&����CU�
NךU���u�u�;���<����&����D��F�����
�0�
�f�g�m�W���H����_��=N��U���u�0�
�b�l�}�Wϸ�&����J)��hZ�����;�
� �l�c�-�W������^��N�������g��#�k�(݁�����9��R�����u�u�u��/��#ݰ�����l ��_�*��"�0�u�&�;�)�ׁ�����9��^��H��r�u�9�0�]�}�W���Y����f(��r����
�
�
�0��n�G�ԜY�ƪ�l��{:��:���c�
� �d�`��F��Y����@��hX�����d�f�%�n�w�}����4����])��hX�����-�
�
�
�"�l�G܁�K���@��[�����6�:�}�;�>�3�Ǯ�+����G9��h��D��
�f�u�u�9�4��������]��[�*ٓ��|�n�u�w�;�(���5�Ԣ�F��1��*���,�0�3�
�g�j����D���F�N�����<�l�6�&��<����&����l��@��U¦�9�!�%�
�d�;�(��H����O�I�\ʰ�&�u�u�u�w�}�������� 9��h_�B���n�u�u�3���;���6����9��Q��Lڊ�f�i�u�u�w�}�Wϸ�&����gT��B��@���
�c�
�d� �8�Wǭ�����9��h[�*��e�u�u�d�~�8����Y���F��Y1�����%�6�0��2��B�ԜY�ƪ�l��{:��:���c�
� �`�o�-�W��	����F
��W�� ���c�%�n�u�w�;�(���5�Ԣ�F��1��*���
�
�
� �c�k����Dӕ��l
��^�����'� �&�2�2�u�(�������l ��V�����~� �&�2�2�u��������EW��G����u��-� ��3����L����U��G�� ��e�%�u�h�]�}�W���Y����9��T��*���!�3�
�`��n� ���Yە��l��1�����b�
�g�e�w�}�F�������9F�N��U���
�8�
�
�"�i�G���B��� ��O#��!ػ� �
�a�d�1��Oׁ�J���9F�N��U���-� ��;�"��C���&����CW��_��]���
�8�m�<�1��O݁�K���F�G�����_�u�u�u�w�3�'�������9��UךU����-� ��9�(�(�������9��R�����&�9�
�d�1��Bہ�L���F��h��9����!�m�
�9�8����H����_��G\��Hʦ�1�9�2�6�!�>��������V��h<�� ���c�
� �g�a�-�^�������]��V�����
�#�m�f���^�ԜY�ƪ�l��{:��:���m�
�;�3��-�(���K�ޓ� F�d��U���u�'�!�g�>�4����
����@��B1�E���u�=�;�}�2���������lT��h�E���u�d�|�0�$�}�W���Y����V
��Z��G���
�`�
�f�]�}�W��Y����U��_��ʴ�&�2�u�'�4�.�Y��s���T��Q��Fۊ�0�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��*���u�%�&�2�4�8�(���
�ғ�@��N��*���
�&�$���)�F���������D�����
��&�d��.�(��Y����Z��D��&���!�f�3�8�f�q����&����|��V�����f�b�u�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����ޓ�@�� B�����2�6�0�
��.�E߁�
����F��h��*���$��
�!�n�;���P�����^ ךU���u�u�3�}�9�)�_�������l
��^��U���%�6�|�u�%�u��������\��h_��U���&�2�6�0��	��������F��F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�8�}��������_	��T1�Hʴ�
�<�
�&�&��(���K����lW����]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�e�}����	����@��X	��*���u�%�&�2�4�8�(���
����U��X�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��@��CN�����:�&�
�:�>��^�������C9��Y�����6�d�h�4��4�(�������@��h��*��u�;�u�4��2����¹��F��X��2��� �
�m�'�0�l�C���Y�����T�����d�e�h�7�8��0�������l��h_�B���;�u�4�
�8�.�(�������F��h��*���$��
�!�n�;���P�ƣ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�l�u�;�w�<�(���
����9��
N������,� �
�o�/���M���F��R ��U���u�u�u�u�0�-����J¹��Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�'�
�"�l�F���Y����C9��Y�����6�d�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z�������lW��h����2�u�'�6�$�s�Z�ԜY�ƫ�C9��h_�*���4�&�2�
�%�>�MϮ�������D�����
��&�d�1�0�G������� J��R	��B���6�
������������V9��1��*��
�f�u�%�$�:����&����GS��D��Yʳ�
���,�"�����	����
9��P1�F���4�
�<�
�$�,�$����ғ�@��B�����2�6�0�
��.�O������R��^	������
�!�m�1�0�F���Y����V��=N��U���u�3�}�4��2��������F�V�����&�$��
�#�e����H���G��d��U���u�u�u�2�'�;�(��&���F��P1�M�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��]��U���;�_�u�u�w�}�W�������lW��h�I����-� ���)�:������� _��R	��F��_�u�u�u�w�1����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�m�3�:�j�^������F�N��U���2�%�3�
�d��G��Y����Q��=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�F��������YNךU���u�u�u�u�%����H����[��[1��0����:�!� ��j����H����_��G]�U���u�u�0�&�w�}�W���Y�����h��D���%�u�h�w���/���!����k>��o6��-������w�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƫ�C9��h_�*��4�&�2�u�%�>���T���F��G1��*��
�d�4�&�0�����CӖ��P�������6�0�
��$�l����I�ƥ�l0��B�����c�y�3�
���#���&����U��\��F���%�&�2�6�2��#���L����lR�Q=��0���� �
�m�1��Aف�J�ƭ�l��h�����
�!�a�3�:�l�[Ͽ�&����P��h=�����3�8�b�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��M���8�d�|�u�?�3�}���Y���F�P�����f�
�d�i�w�-��������9��^�E��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������F9��1��U��3�
����(�(�������9��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���ׁ�
����F��R ��U���u�u�u�u�0�-����J¹��Z�E��D��_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����l ��hZ��U���;�_�u�u�w�}�W�������lW��h�I��������)�F�������9��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���ށ�
����F��R ��U���u�u�u�u�0�-����J¹��Z�^ ����_�u�u�u�w�1��ԜY���F�N�����
�f�
�d�k�}�/���!����k>��o6��-���������L���Y�������U���u�0�1�%�8�8��Զs���K��E�� ��b�%�u�&�>�3�������KǻN����� �d�b�%��.����	����	F��X��¼�
�$�f�u�'�.��������l��h��*���4�
�<�
�$�,�$���ǹ��^9��������;� �
�c�l����H������u;��9���'�
�m�0�e�/���J����C9��P1������&�d�
�$��E�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�f�����K����[��=N��U���u�u�u�'��(�F���	�����u;��9���'�
�m�0�e�/���J��ƹF�N�����u�}�%�6�9�)���������D�����
��&�b�1�0�A�������9F�N��U���u�'�
� �f�j����Dӏ��e��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$���ہ�
����F��R ��U���u�u�u�u�0�-����JĹ��Z�Q=��8���g��!�m������K����F�N�����u�u�u�u�w�}�WϹ�	����U��G^��H���������/���!����k>��o6��-���_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������lW��h�����2�
�'�6�m�-����
ۏ��c*��V��*Ҋ�
�y�<�
��h�W���&������D�����
��&�b�1�0�A���	����l��F1��*���
�&�
�y�6�����
����g9��]�����g�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��Dي�&�
�g�|�#�8�W���Y���F�	��*���d�b�%�u�j�4�(���L���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���2�%�3�
�d��F��Y����*��^ ��M���e�_�u�u�w�}����Y�έ�l��D�����
�u�u�%�$�:����&����GR��D��\���=�;�_�u�w�}�W���Y����U��Y��D��u�0�
�c�l�}�W���YӃ��VFǻN��U���u�u�'�
�"�l�@���Y���k>��o6��-���������/���!����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���2�%�3�
�c�����Ӈ��Z��G�����u�x�u�u�0�-����M����P	��h�����%�:�u�u�%�>����	����l��F1��*���d�3�8�d�{�)���&����U��N�����%�d�<�'�0�l�G��
����^��h�����f�g�u�0��0�Eց�&����U��N�����%�b�<�'�0�l�E������T9��R��!���d�
�&�
�f�}��������B9��h��B���8�d�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���b�3�8�d�~�}����s���F�N�����3�
�a�
�'�2���Y����\��h��*��u�u�u�u�2�.����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\ʴ�1�}�%�6�9�)����I����V
��Z�*���0�
�f�m�w�3�Wǿ�&����G9��1�Hʦ�9�!�%�b�>�/���K����]��X�����:�&�
�#��}�W���&����9��E��D��|�|�u�=�9�W�W���Y���F��G1��*��
�%�:�0�k�}��������ES��d��U���u�0�&�3��u��������\��h_��U���&�2�6�0��	���&����W�V ��]���6�;�!�9�f�m�JϪ�	����A��]�\ʴ�1�}�%�6�9�)����I����V
��Z�*���0�
�f�c�w�3�Wǿ�&����G9��1�Hʦ�9�!�%�e�>�/���H����]�V�����
�#�
�u�w�8�(���Kʹ��A��]�\ʴ�1�}�%�6�9�)����I����V
��Z�*���0�
�f�a�~�}����s���F�N�����3�
�a�
�'�2���Y����\��h��*��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������F9��1�����u�h�4�
�8�.�(���&��ƹF�N�����_�u�u�u�w�}�W���&����U��G����u����l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����A��B1�F���u�&�<�;�'�2����Y��ƹF��E�� ��f�%�
�&�>�3����Y�Ƽ�\��DF��*���'�;�0�l�2�l�W���)����Z��1��D���0�
�b�y�6�����
����g9��_�����e�u�8�
�e�/���I����V
��Z�*���0�
�f�c�w�8�(���Kù��A��]�Yʦ�9�!�%�l�>�/���H����V
��Z�*���0�
�f�a�w�-��������`2��C_�����d�y�4�
�>�����*����Q��D��C�ߊu�u�0�<�]�}�W���Y���N��h�����:�<�
�u�w�-��������`2��C_�����d�|�:�u��-��������Z��S�����2�6�0�
��.�F݁�
����F��SN�����;�!�9�d�g�`��������l��R	��F��u�;�u�4��2����¹��F��[1�����<�'�2�d�e�t�������R��X ��*���
�u�u�0��0�E߁�&����U��G��\ʡ�0�u�u�u�w�}�W�������F9��1��U��'�2�d�m�]�}�W���Y����UF������!�9�2�6�f�`��������V��c1��D؊�&�
�d�u�9�}��������_��N�����`�
�0�
�d�m�W���Yۇ��P	��C1��D��h�&�9�!�'�l��������O��Y
�����:�&�
�#��}�W���&����9��E��D��|�4�1�}�'�>�����ד�[��R����
�
�0�
�d�e�W���Yۇ��P	��C1��D��h�&�9�!�'�j��������O����ߊu�u�u�u�w�}��������l��S������4�;�
���L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�g�t����Y���F�N��U���
� �d�f�'�}�JϷ�&����R��hW��*��u�u�u�u�2�.�W���Y���F�	��*���d�f�%�u�j��/���!����k>��o6��-���������}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��G1��*��
�d�4�&�0�}����
���l�N�����
�a�
�d�6�.���������T��]�����4�2���(������T9��R��!���d�
�&�
�g�}����K����lW��B�����8�d�
�
�2��D��Y����G��1�����d�d�y�&�;�)��������lW��B�����8�f�
�
�2��D��Y����Z��D��&���!�g�3�8�f�q��������V��c1��D݊�&�
�c�_�w�}����s���F�^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�a�t����Y���F�N��U���
� �d�f�'�}�JϿ�&����G9��\��3��e�e�_�u�w�}�W��������T�����2�6�d�h�6�����
����g9��\�����d�u�;�u�6�����&����F�C��@؊�0�
�f�e�w�3�Wǿ�&����G9��1�Hʦ�9�!�%�d�>�/���I����]�V�����
�#�
�u�w�8�(���Kù��A��]�\ʴ�1�}�%�6�9�)����I����V
��Z�*���0�
�f�m�w�3�Wǿ�&����G9��1�Hʦ�9�!�%�b�>�/���K�����YNךU���u�u�u�u�%����J����[��G1�����9�f�
�n�w�}�W�������N�V�����
�:�<�
�w�}��������B9��h��D���8�d�|�:�w�u��������\��h_��U���&�2�6�0��	���&����W�V ��]���6�;�!�9�f�m�Jϭ�����_��h��*��m�u�;�u�6�����&����F�D�����b�<�'�2�f�o�^Ͽ�ӈ��N��h�����#�
�u�u�2����&����T9��\��\���!�0�u�u�w�}�W���YӁ��l ��Z�����h�<�
��%�3��������F�N�����u�u�u�u�w�}�WϹ�	����R��G_��H���������/���!����k>��o6��-���_�u�u�u�w�3�W���Y����������n�_�u�u�9�/����M����W9��V
�� ��
�g�i�u�g�c����
����F��_��H��r�n�u�u�;�>�!��&����W��GZ��Hʥ��9�
�a�1��G���	������Y��G���_�u�u�:���F���&����l��S��*���g�b�
� �f�l�(��K���F��@ ��U���_�u�u�:���(���M�ԓ�F������&�3�
�e��l�E���Y�ƨ�D��^����u�:�
�
��(�E���	��� ��b ��;���!�'�
�g�1��Gف�H����W	��C��F��u�u�9�6��n����Kù��Z�Q=��;�����0�8�e����O����U�_�����:�e�n�u�w�1����M����W��GZ��Hʥ��9�
�e�1��Gց�H����W	��C��F��u�u�9�6��h����K����Z�G1��؊�e�3�
�e��l�E���Y�ƨ�D��^����u�:�
�
��(�A���	�����V��Bۊ� �c�`�%��m��������]ǻN�����
�
� �c�n�-�W��	����9��h��C���%�}�f�x�f�9� ���Y����F�[��#���3�
�m�
�c�a�W����ԓ�9��hX�*��f�u�:�;�8�o�^�ԜY�Ơ�P9��1��*��
�d�i�u��<�E��&����W��F�U���u�:�;�:�g�f�W�������l ��_�����h�%��9�����A���� V��X����|�_�u�u�8�1�ށ�����l��S��E���=�;�}�:���(���O�ӓ�F�V�����
�#�
��w�1����[���F��C��G���
�f�
�g�k�}�G������_	��a1�����a�
�a�h�6�����&����u �R��U��n�u�u�;�#�5�D���&����CT�
N��Wʢ�0�u�9�6��i����H����[��G1�����9�m��|�2�.�W��B�����[��*���l�g�%�u�j��Uϩ�����^��1��*��
�a�h�4��2����˹��F��D��D��u�u�;�!�?����O����[�L�����}�:�
�
��(�E���	���R��X ��*���
��u�9�2��U�ԜY�Ƣ�G��1��*��
�g�i�u�f�}����Q����e9��Q��Lߊ�d�h�4�
�8�.�(���J���V
��L�N���u�;�!�=�e�;�(��&���F�N�����9�6��b�1��Bց�H����C9��Y����
�|�0�&�w�m�L���Yӈ��A��h��B���%�u�h�w�u�*��������lS��B1�F���u�u�%�6�9�)���&����_��^�����u�:�'�&��(�N���	���D�������8�
�d�3��e�(��DӇ��P	��C1��Gي�|�0�&�u�g�f�W���	����9��^1��*��
�f�i�u�w�}�W�������]��[�*���=�;�}�8��l����H����V�
N��R���9�0�_�u�w�}�W���&����U��^��D�ߊu�u�
�a�b�l����Kù��Z�=N��U���u�%�6�;�#�1�E܁�Y����N��G1�*���`�a�%�}�~�`�P���Y����l�N��Uʹ�6��d�3��o�(��s���C9��[��*���d�g�
�f�k�}�W���Y����C9��Y����
�u�=�;��0�(�������W��F�U���d�|�0�&�w�}�W���Yӊ��l0��1��*��l�%�n�u�w�-�%�������l ��[�����h�}�
�4�e�.����I˹��U��S�����d�u�u�8��i����M˹��]ǻN��*��� �!�c�
�"�o�A���Y���R��X ��*���e�e�s�9�4��E���&����CR�=N��U���0� �!�c��(�D���	���N��h;�� ����0�8�g��(�E���	������Y��F���s�!�%�b�����O����l�N��'���9�
�g�3��m�B���Y���R��X ��*���e�e�s�9�4��F߁�����
9��UךU���
�0� �!�a����O����Z������b�
� �d�f��F��Y����G	�G��U���
�b�3�
�f�h����s���C9��D��*��� �a�m�%�w�`�_�������l
��1�Sʹ�6��3�
�f��C��Y����l0��1�*���c�l�%�u�j�/���A���F��a��*���3�
�a�
�f�a�W���)����]��1��E�ߊu�u�
�4�e�j�(���O�ד�F���%���4�2�
�
��f�W���	����9��h��D��
�d�i�u�;��9�������^��h\�����f�e�_�u�w�����
����V��G_��Hʼ�
�'�1�-�2�)��������9F������<�3�
�e��n�K���Y���F��d1��9����!�d�m�%�:�F��Y����N��G1�*���
�f�e�e�w�}�F�������9F�N��U�������#�l�A���&����CU��N�����d�<�l�6�$���������_��N�U���u�u�u�4��2�����ӓ�V��_��]���
�
�d�g��(�F��&���F�_��U���0�_�u�u�w�}��������EW��^����u�0�
�
��<����
����lR��h�I���u�u�u�u�6�����&����lS�������8�
�
�
�c�;�(��&���F�_��U���0�_�u�u�w�}��������EW��^����u�0�
�
���(�������G9��h\�*��i�u�u�u�w�}��������_��h[�U���;�}�8�
���(�������9��^��H��r�u�9�0�]�}�W���Y����\��h��@��e�_�u�u�2��F���&����l��S��U���u�u�4�
�8�.�(���L����F��R �����<�<�
�b�1��G���	����[�I�����u�u�u�u�w�<�(���
����S��^����u�0�
�
�"�i�O���Y���F�N�����:�&�
�#�b�i�G������G��^1��Gފ� �a�g�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�B��I��ƹF��R��*���
� �g�c�'�}�J�ԜY���F��h�����#�`�a�e�w�5��������Z9��[�� ��e�%�}�|�j�z�P������F�N�����:�&�
�#�b�i�G��Y����V
��Z�*��� �m�l�%�w�`�_���&����U��N��U���
�e�
�0�8�:��������
9��UךU���0�
�8�d����������l��S�����!�%�d�<�1��Fց�KӞ����T�����d�d�n�u�w�.����	�ԓ�l ��_�����h�_�u�u�w�}�$���5����F��V�����g�g�"�0�w�.����	�ד�l��h_�C��u�u�d�|�2�.�W���Y�����C�����
�e�
�f�]�}�W���&����9��S�����
� �m�`�'�}�J�������l �� [�����'�&�9�!�'�l����&����CT�=N��U���
�8�d�
��(�O���	���N��[1�����<�1�8�'�6����L����K	��V�����
�#�
�|�]�}�W���&����
9��Q��F݊�g�i�u�!�'�i�(���N�ߓ�F��EN��*���&�
�#�
�~�W�W�������CW��B1�M���u�h�w�w� �8�WǸ�&����gT��B��@���
�%�,�0�1��O߁�J����C9��Y����
�e�|�0�$�}�G��Y����V
��Z��؊� �g�c�%�w�`�_���&����Z9��h\�*��-�'�4�
�8�.�(���&����F�D�����
�f�3�
�g�h����D�θ�C9��^_�� ��f�
�g�-�%�<�(���
����9��d��Uʦ�9�!�%�
��(�C���	���N��G1�����
�g�
�g�/�/��������_��G�U���&�9�!�%�g�4����M����Z���*���d�
�
� �o�l�����ƿ�_9��G_�����
�f�
�g�l�}�Wϭ�����W��h��L���%�u�h�_�w�}�W���*����v%��B��AҊ�0�
�g�g� �8�Wǭ�����V��h��*��g�e�u�u�f�t����Y���F���*���d�
�
� �n�m���Y����V
��Z�*��� �m�`�%�w�`�_���&�ד�F9��1��U���u�0�
�8�f��(���&����_��G�U���&�9�!�%�n�4����O¹��Z���*���3�
�e�
�e�<�ϭ�����^��h��M���%�|�_�u�w�8�(���K����^��G\��H���0�
�8�
�"�h�E���Y����V
��Z�����b�
�g�n�w�}��������ZT��B1�G���u�h�}�8��n�(���&����lT��h����&�9�!�%��o����OŹ��]ǻN�����8�g�<�
�"�l�Oށ�K�����h_�*���d�3�
�e�d�-�W���Y����G��h�����e�`�%�|�]�}�W���&����l��B1�A���u�h�}�8��n�(���&����P��N��ʦ�9�!�%�
��(�C���	����F�D�����e�<�3�
�e��D��Y���F���&�����!�d�o�/���N�ƻ�V�D�����l�<�'�2�f�l�_���D����F��D��U���u�u�&�9�#�-�F�������9��d��Uʦ�9�!�%�b�>�;�(��&���F��Z��@���
�m�
�g�6�9��������l��B1�D���|�_�u�u�2����&����l_��h�I���u�u�u�u�6�����&����lQ��^�Eʢ�0�u�&�9�#�-�F������� V��G��U��|�0�&�u�w�}�W�������A��^��G���
�l�
�f�]�}�W���&����9��Q��Aۊ�f�i�u�u�w�}�Wϸ�&����9��1�����l�
�f�"�2�}��������l��R	��F��e�u�u�d�~�8����Y���F��R����
�
� �l�c�-�L���Yӕ��l��W��*���l�m�%�u�j�W�W���Y�ƥ�l6��E�����0�e�"�0�w�.����	�ߓ�l��h_�M��u�u�d�|�2�.�W���Y�����h��@ڊ�
� �l�d�'�f�W���
����^��Q��D���%�u�h�w�u�*��������f*��Y!��*���<�
�%�,�2�;�(��N����F��h�����#�`�a�e�~�8����I��ƹF��R�����<�3�
�b��o�K���H�ƻ�V�Q=��8���g��!�m��3����	����lT��h�Hʴ�
�:�&�
�!�h�C��PӃ��VF�UךU���0�
�8�b�1��F���	���D��������-� ��9�(�(�������g��h��D��
�f�h�4��2�����ӓ�V�R��U��n�u�u�&�;�)�؁�&����P��N�U��u�=�;�}��%�"�������R��Y1��!���
� �g�m�'�}�W�������l
��1�E���9�0�w�w�]�}�W���&����l ��_�*��i�u�&�9�#�-�(���H����CT��EN�����%�
� �d�o��E��Y����V
��Z�����
�m�
�g�k�}��������Z9��h]�*��:�u�0�
�:�j����&����CT�=N��U���
�8�
� �b�o����D������YN��&��� ��;� ��h����	����l ��V�����u�%�6�;�#�1�Fځ�M���V
��L�N���u�&�9�!�'�4�(���K�ޓ� F�d��U���u�'�!�<�>�4����JŹ����YN�����
�
�
� �e�i����P���A�R��U���u�u�u�4��2�����ӓ�V��N�����!�%�<�
�"�l�A؁�J���9F�N��U���
�d�3�
�g�h�������G��^1��*���d�f�
�g�g�}�W��PӃ��VFǻN��U���%�6�;�!�;�l�(��B�����h��*��� �a�e�%�w�`�}���Y���A��^1��*��
�f�"�0�w�)��������T��G\��\��r�r�u�9�2�W�W���Y�ƭ�l��D�����a�e�_�u�w�0�(��&����lU��h�I���d�u�=�;��4��������f*��Y!��*���<�
�-�
�����M����Z��^	��´�
�:�&�
�!�e�F�������V�=N��U���
�e�
�0�8�:��������
9��R��]���
�
�f�<�1��E؁�KӇ����h��A���3�
�f�
�e�f�W�������_��R�����<�3�
�b��o�K�������l��^1��*��
�g�4�1�#�-����&����lP��h�N���u�!�%�d�f�9��������U��_��G��u�!�%�<�>��(�������
9����U���
�
�g�<�1��Gځ�K��ƹF��Z��Fۊ�
�d�3�
�g�n����D������YN�����
�e�3�
�g�d����Y����\��h��*���u�9�0�w�u�W�W�������9��^1��*��
�g�i�u�f�}����Q����e9��hZ�*��h�4�
�:�$��ׁ�?�Ʃ�@�L�U���!�%�d�d�>�4����&����CT�
N��Wʢ�0�u�9�6��o����Hù��[��G1�����9�m��|�2�.�W��B�����h\�����e�
�g�i�w�l�W����ο�T��������;� �
�b�4�(���&����U��X��G���u�<�;�1�6�����&����lW������w�_�u�u�:��C���&����CU�
N�����e�3�
�a��n�QϮ�I����9��h[�*��n�u�u�!�'�o�(���H����CT�
N��Wʢ�0�u�&�2�2�u�$���,����|��\�����%��d�3��l�D���P����Z��SF��*���&�
�#�m��t�W�������l�N����
� �d�d��o�K���H�ƻ�V�D������-� ��9�(�(�������C9��1��*��f�%�|�i�$�:����	����@��A_��D���0�&�u�e�l�}�WϪ�	����U��[�����h�}�8�
�b�;�(��N����F��Z�*ۊ� �d�g�
�d�f�W�������9��h[�*��i�u�!�%�$�;�(��&����AF��G1�*���`�m�%�|�]�}�W���&�ߓ�F9��1��U��_�u�u�u�w�-��������l ��@��U¡�%�&�3�
�g��E��Y���O��[�����u�u�u�%�4�3����A����F�C��Fڊ� �`�e�%�w�`�}���Y���G��W�� ���m�%�u�=�9�u����A����W��G\��\��r�r�u�9�2�W�W���Y�Ƹ�C9��h��@���%�n�u�u�#�-�Dށ�����l��S�����<�3�
�e��o��������9��Q��E܊�g�n�u�u�#�-�D݁�����l��S��U���u�u�4�
�8�.�(���&����[����*��� �f�e�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�(��Y����^��1��*��
�f�i�u�w�}�W�������9��h]�*��"�0�u�!�'�n�(���J�ԓ�N��S��D���0�&�u�u�w�}�WϪ�	����U��Z��D�ߊu�u�8�
�c�;�(��&���F��Z��*���
�`�3�
�d��Eϱ�Y����[��B1�C���|�_�u�u�:��A���&����CT�
N�����a�'�2�d�a�}��������lW��h�N���u�!�%�f��(�@���	���N��C��D���
�g�
�g�8�}����
¹��lQ��h�N���u�!�%�f��(�@���	���N��C��G���
�a�
�g�8�}����
����lQ��h�N���u�!�%�f��(�@���	���N��G1�*���b�l�%�u�9�}����A����R��G\����u�8�
�d�1��Bց�K�����h]�����`�
�g�4�3�:����&����CT�=N��U���
�g�3�
�`��E��Yۈ��A��h��B���%�u�'�;�#�5�D���&����CT�=N��U���
�f�3�
�o��E��Yے��lR��Q��B݊�g�4�1�!�'�n�(���N�ߓ�O��N�����a�
� �d�n�2����Y����C9��Y�����g�_�u�u�:��C���&����CV�
N����m�_�u�u�:��C���&����CW�
N��*���'�;�0�l�2�l�}���Y����S��B1�L���u�h�}�8��n����A��������*���3�
�a�
�e�f�W�������9��hY�*��i�u�!�%�c����N����R��C��FҊ� �b�b�%�~�W�W�������l ��[�����1�u�h�4��2����ƹ��9F���*���3�
�`�
�g�a�W���&����9F���*���3�
�`�
�f�a�W���)����]��1��E�ߊu�u�8�
�o�;�(��&���F��Z��C���
�l�
�g�6�9����MĹ��lW��h�N���u�!�%�`��(�O���	���N��G1�*���
�g�`�4�3�:����&����CT�=N��U���
�d�3�
�b��������R��X ��*���
�n�u�u�#�-�Bށ�����l��S�����b�n�u�u�#�-�Bށ�����l��S������4�2�
���L���YӒ��lS��Q��E݊�g�i�u�!�'�i�(���N�Փ�F��SN�����
� �d�l�'�t�}���Y����U��B1�Gۊ�g�i�u�!�'�o�(���H����CT��EN����
� �d�d��o�L���YӒ��lS��Q��D���%�u�h�_�w�}�W���	����@��AV��3ʢ�0�u�!�%�e����Iʹ��V�
N��R���9�0�_�u�w�}�W�������l
��h^�U���!�%�`�
�"�l�C؁�J���9F�N��U���
�a�3�
�f�h�������G��]�� ��g�
�g�e�w�}�F�������9F�N��U���
�e�3�
�f�n���Y����^��1��*��
�a�i�u��%�3�������l��^ �����b�
�d�f�w�2����K����F�C��@݊� �d�e�
�e�a�Wǰ�����l ��W�����'�;�!�=�c�;�(��&���9F���*���<�3�
�a��n�K������� 9��h]�*��s�%�e�g���(���J�ޓ� O��N�����m�
� �`�a�-�W������f*��Y!��*���<�
�-�
�����O����F�N�����u�|�_�u�w�0�(�������9��R�������g��#�e�(�������lW��B1�A���}�u�u�u�8�3���B�����hW�����d�f�%�u�j�;�(���5�Ԣ�F��1��*���
�
�
� �f�m�(��A�����Y��E��u�u�!�%�n����A����[��d1��1��� �
�g�!��3�(���@�ғ�N��C��U���;�:�e�n�w�}�������� 9��R��]���
�e�
�0�8�:��������9�������d�d�1�8�%�<�(�������l��d��Uʡ�%�<�3�
�g��E��Y���D��F�����}��-� ��3����M����V��a1�����l�
�g�u�w�4��������]��[�*���|�0�&�u�g�f�W�������l��Y�� ��f�
�g�i�w�l�W����Π�P9��_�� ��g�
�d�h�6�����&����lV�R��U��n�u�u�!�'�4�ށ����� 9��R��W���"�0�u�9�4��F߁�����
9��S�����;�!�9�m�g�}����[����F�C�����
�
�c�3��d�(��E���F��R ������m�3�
�o��C������]��[��3���0�&�u�e�l�}�WϪ�	����9��Q��Cӊ�g�i�u�e�w�5��������9��hX�*��h�4�
�:�$�����I�Ʃ�@�L�U���!�%�<�<�����L����[�L�����}�:�
�
��(�A���	���R��X ��*���f�e�u�9�2��U�ԜY�Ƹ�C9��^]��*���c�b�%�u�j��Uϩ�����\��hZ�� ��f�%�u�u�'�>�����ޓ�uO��[��W���_�u�u�8���C������� 9��R��W���"�0�u�9�4��B���&����CW������!�9�g�
�~�8����H��ƹF��Z��*���<�3�
�c��o�K���H�ƻ�V�[��#���3�
�a�
�c�`��������_��q(�����u�e�n�u�w�)��������U��\��G��u�d�u�=�9�u����&¹��lR��h�Hʴ�
�:�&�
�!�n�G������D��N�����<�<�3�
�e��E��Y���D��F�����3�
�d�
�c�`��������_��G�����w�w�_�u�w�0�(���&����l ��]�����h�w�w�"�2�}����/�Փ�F9��1��U���%�6�;�!�;�o�(�������V�=N��U���
�
�
�
�"�o�C���Y���D��_��]���
�
�
� �e�m����Y����\��h��*���0�&�u�e�l�}�WϪ�	����F9��1��U��w�w�"�0�w�.����Q����~3�� ����
�;�0�%��l����@Ź��F�D�����%�6�;�!�;�l�(���PӃ��VF�U�����0�4�n�